`timescale 1 ns / 1 ns

module simulink_functio_tb;

  reg  clk;
  reg  reset_x;
  wire clk_enable;
  wire alpha_arctangen_done;  // ufix1
  wire rdEnb;
  wire alpha_arctangen_done_enb;  // ufix1
  reg [9:0] magnitude_addr;  // ufix10
  wire alpha_arctangen_lastAddr;  // ufix1
  wire resetn;
  reg  check2_done;  // ufix1
  wire magnitude_done;  // ufix1
  wire magnitude_done_enb;  // ufix1
  wire magnitude_active;  // ufix1
  reg [9:0] Data_Type_Conversion1_out1_addr;  // ufix10
  wire [15:0] in_im_table_data [0:1000];  // ufix16 [1001]
  wire [15:0] in_im_1;  // ufix16
  wire signed [15:0] rawData_in_im;  // sfix16_En14
  reg signed [15:0] holdData_in_im;  // sfix16_En14
  reg signed [15:0] in_im_offset;  // sfix16_En14
  wire signed [15:0] in_im_2;  // sfix16_En14
  wire Data_Type_Conversion1_out1_active;  // ufix1
  reg  tb_enb_delay;
  wire Data_Type_Conversion1_out1_enb;  // ufix1
  wire [15:0] in_re_table_data [0:1000];  // ufix16 [1001]
  wire [15:0] in_re_1;  // ufix16
  wire signed [15:0] rawData_in_re;  // sfix16_En14
  reg signed [15:0] holdData_in_re;  // sfix16_En14
  reg signed [15:0] in_re_offset;  // sfix16_En14
  wire signed [15:0] in_re_2;  // sfix16_En14
  wire snkDone;
  wire snkDonen;
  wire tb_enb;
  wire [15:0] magnitude;  // ufix16_En14
  wire signed [7:0] alpha_arctangen;  // sfix8_En5
  wire magnitude_enb;  // ufix1
  wire magnitude_lastAddr;  // ufix1
  reg  check1_done;  // ufix1
  wire [15:0] magnitude_expected_table_data [0:1000];  // ufix16 [1001]
  wire [15:0] magnitude_expected_1;  // ufix16
  wire [15:0] magnitude_expected_2;  // ufix16_En14
  wire [15:0] magnitude_ref;  // ufix16_En14
  reg  magnitude_testFailure;  // ufix1
  wire [7:0] alpha_arctangen_expected_table_data [0:1000];  // ufix8 [1001]
  wire [7:0] alpha_arctangen_expected_1;  // ufix8
  wire signed [7:0] alpha_arctangen_expected_2;  // sfix8_En5
  wire signed [7:0] alpha_arctangen_ref;  // sfix8_En5
  reg  alpha_arctangen_testFailure;  // ufix1
  wire testFailure;  // ufix1


  assign alpha_arctangen_done_enb = alpha_arctangen_done & rdEnb;



  assign alpha_arctangen_lastAddr = magnitude_addr >= 10'b1111101000;



  assign alpha_arctangen_done = alpha_arctangen_lastAddr & resetn;



  // Delay to allow last sim cycle to complete
  always @(posedge clk)
    begin : checkDone_2
      if (reset_x) begin
        check2_done <= 0;
      end
      else begin
        if (alpha_arctangen_done_enb) begin
          check2_done <= alpha_arctangen_done;
        end
      end
    end

  assign magnitude_done_enb = magnitude_done & rdEnb;



  assign magnitude_active = magnitude_addr != 10'b1111101000;



  // Data source for in_im
  assign in_im_table_data[0] = 16'b1111111111111111;
  assign in_im_table_data[1] = 16'b0000100111010100;
  assign in_im_table_data[2] = 16'b0001010011001100;
  assign in_im_table_data[3] = 16'b0001110111110100;
  assign in_im_table_data[4] = 16'b0010011100011010;
  assign in_im_table_data[5] = 16'b0010111101011000;
  assign in_im_table_data[6] = 16'b0011011011111111;
  assign in_im_table_data[7] = 16'b0011110111100111;
  assign in_im_table_data[8] = 16'b0100001011110110;
  assign in_im_table_data[9] = 16'b0100011111010011;
  assign in_im_table_data[10] = 16'b0100110001100001;
  assign in_im_table_data[11] = 16'b0100110011110010;
  assign in_im_table_data[12] = 16'b0100111101011000;
  assign in_im_table_data[13] = 16'b0100111101011000;
  assign in_im_table_data[14] = 16'b0100110011110010;
  assign in_im_table_data[15] = 16'b0100110001100001;
  assign in_im_table_data[16] = 16'b0100011111010011;
  assign in_im_table_data[17] = 16'b0100001011110110;
  assign in_im_table_data[18] = 16'b0011110111100111;
  assign in_im_table_data[19] = 16'b0011011011111111;
  assign in_im_table_data[20] = 16'b0010111101011000;
  assign in_im_table_data[21] = 16'b0010011100011010;
  assign in_im_table_data[22] = 16'b0001110111110100;
  assign in_im_table_data[23] = 16'b0001010011001100;
  assign in_im_table_data[24] = 16'b0000100111010100;
  assign in_im_table_data[25] = 16'b1111111111111111;
  assign in_im_table_data[26] = 16'b1111011000101011;
  assign in_im_table_data[27] = 16'b1110101100110011;
  assign in_im_table_data[28] = 16'b1110001000001011;
  assign in_im_table_data[29] = 16'b1101100011100101;
  assign in_im_table_data[30] = 16'b1101000010100111;
  assign in_im_table_data[31] = 16'b1100100100000000;
  assign in_im_table_data[32] = 16'b1100001000011000;
  assign in_im_table_data[33] = 16'b1011110100001001;
  assign in_im_table_data[34] = 16'b1011100000101100;
  assign in_im_table_data[35] = 16'b1011001110011110;
  assign in_im_table_data[36] = 16'b1011001100001101;
  assign in_im_table_data[37] = 16'b1011000010100111;
  assign in_im_table_data[38] = 16'b1011000010100111;
  assign in_im_table_data[39] = 16'b1011001100001101;
  assign in_im_table_data[40] = 16'b1011001110011110;
  assign in_im_table_data[41] = 16'b1011100000101100;
  assign in_im_table_data[42] = 16'b1011110100001001;
  assign in_im_table_data[43] = 16'b1100001000011000;
  assign in_im_table_data[44] = 16'b1100100100000000;
  assign in_im_table_data[45] = 16'b1101000010100111;
  assign in_im_table_data[46] = 16'b1101100011100101;
  assign in_im_table_data[47] = 16'b1110001000001011;
  assign in_im_table_data[48] = 16'b1110101100110011;
  assign in_im_table_data[49] = 16'b1111011000101011;
  assign in_im_table_data[50] = 16'b1111111111111111;
  assign in_im_table_data[51] = 16'b0000100111010100;
  assign in_im_table_data[52] = 16'b0001010011001100;
  assign in_im_table_data[53] = 16'b0001110111110100;
  assign in_im_table_data[54] = 16'b0010011100011010;
  assign in_im_table_data[55] = 16'b0010111101011000;
  assign in_im_table_data[56] = 16'b0011011011111111;
  assign in_im_table_data[57] = 16'b0011110111100111;
  assign in_im_table_data[58] = 16'b0100001011110110;
  assign in_im_table_data[59] = 16'b0100011111010011;
  assign in_im_table_data[60] = 16'b0100110001100001;
  assign in_im_table_data[61] = 16'b0100110011110010;
  assign in_im_table_data[62] = 16'b0100111101011000;
  assign in_im_table_data[63] = 16'b0100111101011000;
  assign in_im_table_data[64] = 16'b0100110011110010;
  assign in_im_table_data[65] = 16'b0100110001100001;
  assign in_im_table_data[66] = 16'b0100011111010011;
  assign in_im_table_data[67] = 16'b0100001011110110;
  assign in_im_table_data[68] = 16'b0011110111100111;
  assign in_im_table_data[69] = 16'b0011011011111111;
  assign in_im_table_data[70] = 16'b0010111101011000;
  assign in_im_table_data[71] = 16'b0010011100011010;
  assign in_im_table_data[72] = 16'b0001110111110100;
  assign in_im_table_data[73] = 16'b0001010011001100;
  assign in_im_table_data[74] = 16'b0000100111010100;
  assign in_im_table_data[75] = 16'b1111111111111111;
  assign in_im_table_data[76] = 16'b1111011000101011;
  assign in_im_table_data[77] = 16'b1110101100110011;
  assign in_im_table_data[78] = 16'b1110001000001011;
  assign in_im_table_data[79] = 16'b1101100011100101;
  assign in_im_table_data[80] = 16'b1101000010100111;
  assign in_im_table_data[81] = 16'b1100100100000000;
  assign in_im_table_data[82] = 16'b1100001000011000;
  assign in_im_table_data[83] = 16'b1011110100001001;
  assign in_im_table_data[84] = 16'b1011100000101100;
  assign in_im_table_data[85] = 16'b1011001110011110;
  assign in_im_table_data[86] = 16'b1011001100001101;
  assign in_im_table_data[87] = 16'b1011000010100111;
  assign in_im_table_data[88] = 16'b1011000010100111;
  assign in_im_table_data[89] = 16'b1011001100001101;
  assign in_im_table_data[90] = 16'b1011001110011110;
  assign in_im_table_data[91] = 16'b1011100000101100;
  assign in_im_table_data[92] = 16'b1011110100001001;
  assign in_im_table_data[93] = 16'b1100001000011000;
  assign in_im_table_data[94] = 16'b1100100100000000;
  assign in_im_table_data[95] = 16'b1101000010100111;
  assign in_im_table_data[96] = 16'b1101100011100101;
  assign in_im_table_data[97] = 16'b1110001000001011;
  assign in_im_table_data[98] = 16'b1110101100110011;
  assign in_im_table_data[99] = 16'b1111011000101011;
  assign in_im_table_data[100] = 16'b1111111111111111;
  assign in_im_table_data[101] = 16'b0000100111010100;
  assign in_im_table_data[102] = 16'b0001010011001100;
  assign in_im_table_data[103] = 16'b0001110111110100;
  assign in_im_table_data[104] = 16'b0010011100011010;
  assign in_im_table_data[105] = 16'b0010111101011000;
  assign in_im_table_data[106] = 16'b0011011011111111;
  assign in_im_table_data[107] = 16'b0011110111100111;
  assign in_im_table_data[108] = 16'b0100001011110110;
  assign in_im_table_data[109] = 16'b0100011111010011;
  assign in_im_table_data[110] = 16'b0100110001100001;
  assign in_im_table_data[111] = 16'b0100110011110010;
  assign in_im_table_data[112] = 16'b0100111101011000;
  assign in_im_table_data[113] = 16'b0100111101011000;
  assign in_im_table_data[114] = 16'b0100110011110010;
  assign in_im_table_data[115] = 16'b0100110001100001;
  assign in_im_table_data[116] = 16'b0100011111010011;
  assign in_im_table_data[117] = 16'b0100001011110110;
  assign in_im_table_data[118] = 16'b0011110111100111;
  assign in_im_table_data[119] = 16'b0011011011111111;
  assign in_im_table_data[120] = 16'b0010111101011000;
  assign in_im_table_data[121] = 16'b0010011100011010;
  assign in_im_table_data[122] = 16'b0001110111110100;
  assign in_im_table_data[123] = 16'b0001010011001100;
  assign in_im_table_data[124] = 16'b0000100111010100;
  assign in_im_table_data[125] = 16'b1111111111111111;
  assign in_im_table_data[126] = 16'b1111011000101011;
  assign in_im_table_data[127] = 16'b1110101100110011;
  assign in_im_table_data[128] = 16'b1110001000001011;
  assign in_im_table_data[129] = 16'b1101100011100101;
  assign in_im_table_data[130] = 16'b1101000010100111;
  assign in_im_table_data[131] = 16'b1100100100000000;
  assign in_im_table_data[132] = 16'b1100001000011000;
  assign in_im_table_data[133] = 16'b1011110100001001;
  assign in_im_table_data[134] = 16'b1011100000101100;
  assign in_im_table_data[135] = 16'b1011001110011110;
  assign in_im_table_data[136] = 16'b1011001100001101;
  assign in_im_table_data[137] = 16'b1011000010100111;
  assign in_im_table_data[138] = 16'b1011000010100111;
  assign in_im_table_data[139] = 16'b1011001100001101;
  assign in_im_table_data[140] = 16'b1011001110011110;
  assign in_im_table_data[141] = 16'b1011100000101100;
  assign in_im_table_data[142] = 16'b1011110100001001;
  assign in_im_table_data[143] = 16'b1100001000011000;
  assign in_im_table_data[144] = 16'b1100100100000000;
  assign in_im_table_data[145] = 16'b1101000010100111;
  assign in_im_table_data[146] = 16'b1101100011100101;
  assign in_im_table_data[147] = 16'b1110001000001011;
  assign in_im_table_data[148] = 16'b1110101100110011;
  assign in_im_table_data[149] = 16'b1111011000101011;
  assign in_im_table_data[150] = 16'b1111111111111111;
  assign in_im_table_data[151] = 16'b0000100111010100;
  assign in_im_table_data[152] = 16'b0001010011001100;
  assign in_im_table_data[153] = 16'b0001110111110100;
  assign in_im_table_data[154] = 16'b0010011100011010;
  assign in_im_table_data[155] = 16'b0010111101011000;
  assign in_im_table_data[156] = 16'b0011011011111111;
  assign in_im_table_data[157] = 16'b0011110111100111;
  assign in_im_table_data[158] = 16'b0100001011110110;
  assign in_im_table_data[159] = 16'b0100011111010011;
  assign in_im_table_data[160] = 16'b0100110001100001;
  assign in_im_table_data[161] = 16'b0100110011110010;
  assign in_im_table_data[162] = 16'b0100111101011000;
  assign in_im_table_data[163] = 16'b0100111101011000;
  assign in_im_table_data[164] = 16'b0100110011110010;
  assign in_im_table_data[165] = 16'b0100110001100001;
  assign in_im_table_data[166] = 16'b0100011111010011;
  assign in_im_table_data[167] = 16'b0100001011110110;
  assign in_im_table_data[168] = 16'b0011110111100111;
  assign in_im_table_data[169] = 16'b0011011011111111;
  assign in_im_table_data[170] = 16'b0010111101011000;
  assign in_im_table_data[171] = 16'b0010011100011010;
  assign in_im_table_data[172] = 16'b0001110111110100;
  assign in_im_table_data[173] = 16'b0001010011001100;
  assign in_im_table_data[174] = 16'b0000100111010100;
  assign in_im_table_data[175] = 16'b1111111111111111;
  assign in_im_table_data[176] = 16'b1111011000101011;
  assign in_im_table_data[177] = 16'b1110101100110011;
  assign in_im_table_data[178] = 16'b1110001000001011;
  assign in_im_table_data[179] = 16'b1101100011100101;
  assign in_im_table_data[180] = 16'b1101000010100111;
  assign in_im_table_data[181] = 16'b1100100100000000;
  assign in_im_table_data[182] = 16'b1100001000011000;
  assign in_im_table_data[183] = 16'b1011110100001001;
  assign in_im_table_data[184] = 16'b1011100000101100;
  assign in_im_table_data[185] = 16'b1011001110011110;
  assign in_im_table_data[186] = 16'b1011001100001101;
  assign in_im_table_data[187] = 16'b1011000010100111;
  assign in_im_table_data[188] = 16'b1011000010100111;
  assign in_im_table_data[189] = 16'b1011001100001101;
  assign in_im_table_data[190] = 16'b1011001110011110;
  assign in_im_table_data[191] = 16'b1011100000101100;
  assign in_im_table_data[192] = 16'b1011110100001001;
  assign in_im_table_data[193] = 16'b1100001000011000;
  assign in_im_table_data[194] = 16'b1100100100000000;
  assign in_im_table_data[195] = 16'b1101000010100111;
  assign in_im_table_data[196] = 16'b1101100011100101;
  assign in_im_table_data[197] = 16'b1110001000001011;
  assign in_im_table_data[198] = 16'b1110101100110011;
  assign in_im_table_data[199] = 16'b1111011000101011;
  assign in_im_table_data[200] = 16'b1111111111111111;
  assign in_im_table_data[201] = 16'b0000100111010100;
  assign in_im_table_data[202] = 16'b0001010011001100;
  assign in_im_table_data[203] = 16'b0001110111110100;
  assign in_im_table_data[204] = 16'b0010011100011010;
  assign in_im_table_data[205] = 16'b0010111101011000;
  assign in_im_table_data[206] = 16'b0011011011111111;
  assign in_im_table_data[207] = 16'b0011110111100111;
  assign in_im_table_data[208] = 16'b0100001011110110;
  assign in_im_table_data[209] = 16'b0100011111010011;
  assign in_im_table_data[210] = 16'b0100110001100001;
  assign in_im_table_data[211] = 16'b0100110011110010;
  assign in_im_table_data[212] = 16'b0100111101011000;
  assign in_im_table_data[213] = 16'b0100111101011000;
  assign in_im_table_data[214] = 16'b0100110011110010;
  assign in_im_table_data[215] = 16'b0100110001100001;
  assign in_im_table_data[216] = 16'b0100011111010011;
  assign in_im_table_data[217] = 16'b0100001011110110;
  assign in_im_table_data[218] = 16'b0011110111100111;
  assign in_im_table_data[219] = 16'b0011011011111111;
  assign in_im_table_data[220] = 16'b0010111101011000;
  assign in_im_table_data[221] = 16'b0010011100011010;
  assign in_im_table_data[222] = 16'b0001110111110100;
  assign in_im_table_data[223] = 16'b0001010011001100;
  assign in_im_table_data[224] = 16'b0000100111010100;
  assign in_im_table_data[225] = 16'b1111111111111111;
  assign in_im_table_data[226] = 16'b1111011000101011;
  assign in_im_table_data[227] = 16'b1110101100110011;
  assign in_im_table_data[228] = 16'b1110001000001011;
  assign in_im_table_data[229] = 16'b1101100011100101;
  assign in_im_table_data[230] = 16'b1101000010100111;
  assign in_im_table_data[231] = 16'b1100100100000000;
  assign in_im_table_data[232] = 16'b1100001000011000;
  assign in_im_table_data[233] = 16'b1011110100001001;
  assign in_im_table_data[234] = 16'b1011100000101100;
  assign in_im_table_data[235] = 16'b1011001110011110;
  assign in_im_table_data[236] = 16'b1011001100001101;
  assign in_im_table_data[237] = 16'b1011000010100111;
  assign in_im_table_data[238] = 16'b1011000010100111;
  assign in_im_table_data[239] = 16'b1011001100001101;
  assign in_im_table_data[240] = 16'b1011001110011110;
  assign in_im_table_data[241] = 16'b1011100000101100;
  assign in_im_table_data[242] = 16'b1011110100001001;
  assign in_im_table_data[243] = 16'b1100001000011000;
  assign in_im_table_data[244] = 16'b1100100100000000;
  assign in_im_table_data[245] = 16'b1101000010100111;
  assign in_im_table_data[246] = 16'b1101100011100101;
  assign in_im_table_data[247] = 16'b1110001000001011;
  assign in_im_table_data[248] = 16'b1110101100110011;
  assign in_im_table_data[249] = 16'b1111011000101011;
  assign in_im_table_data[250] = 16'b0000000000000000;
  assign in_im_table_data[251] = 16'b1111110000101001;
  assign in_im_table_data[252] = 16'b1111100100010010;
  assign in_im_table_data[253] = 16'b1111011011011000;
  assign in_im_table_data[254] = 16'b1111001011000001;
  assign in_im_table_data[255] = 16'b1111000100110111;
  assign in_im_table_data[256] = 16'b1110111001011101;
  assign in_im_table_data[257] = 16'b1110110101001101;
  assign in_im_table_data[258] = 16'b1110100111110100;
  assign in_im_table_data[259] = 16'b1110100101001000;
  assign in_im_table_data[260] = 16'b1110011111010011;
  assign in_im_table_data[261] = 16'b1110011110000000;
  assign in_im_table_data[262] = 16'b1110011100001101;
  assign in_im_table_data[263] = 16'b1110011100001101;
  assign in_im_table_data[264] = 16'b1110011110000000;
  assign in_im_table_data[265] = 16'b1110011111010011;
  assign in_im_table_data[266] = 16'b1110100101001000;
  assign in_im_table_data[267] = 16'b1110100111110100;
  assign in_im_table_data[268] = 16'b1110110101001101;
  assign in_im_table_data[269] = 16'b1110111001011101;
  assign in_im_table_data[270] = 16'b1111000100110111;
  assign in_im_table_data[271] = 16'b1111001011000001;
  assign in_im_table_data[272] = 16'b1111011011011000;
  assign in_im_table_data[273] = 16'b1111100100010010;
  assign in_im_table_data[274] = 16'b1111110000101001;
  assign in_im_table_data[275] = 16'b0000000000000000;
  assign in_im_table_data[276] = 16'b0000001111010110;
  assign in_im_table_data[277] = 16'b0000011011101101;
  assign in_im_table_data[278] = 16'b0000100100100111;
  assign in_im_table_data[279] = 16'b0000110100111110;
  assign in_im_table_data[280] = 16'b0000111011001000;
  assign in_im_table_data[281] = 16'b0001000110100010;
  assign in_im_table_data[282] = 16'b0001001010110010;
  assign in_im_table_data[283] = 16'b0001011000001011;
  assign in_im_table_data[284] = 16'b0001011010110111;
  assign in_im_table_data[285] = 16'b0001100000101100;
  assign in_im_table_data[286] = 16'b0001100001111111;
  assign in_im_table_data[287] = 16'b0001100011110010;
  assign in_im_table_data[288] = 16'b0001100011110010;
  assign in_im_table_data[289] = 16'b0001100001111111;
  assign in_im_table_data[290] = 16'b0001100000101100;
  assign in_im_table_data[291] = 16'b0001011010110111;
  assign in_im_table_data[292] = 16'b0001011000001011;
  assign in_im_table_data[293] = 16'b0001001010110010;
  assign in_im_table_data[294] = 16'b0001000110100010;
  assign in_im_table_data[295] = 16'b0000111011001000;
  assign in_im_table_data[296] = 16'b0000110100111110;
  assign in_im_table_data[297] = 16'b0000100100100111;
  assign in_im_table_data[298] = 16'b0000011011101101;
  assign in_im_table_data[299] = 16'b0000001111010110;
  assign in_im_table_data[300] = 16'b0000000000000000;
  assign in_im_table_data[301] = 16'b1111110000101001;
  assign in_im_table_data[302] = 16'b1111100100010010;
  assign in_im_table_data[303] = 16'b1111011011011000;
  assign in_im_table_data[304] = 16'b1111001011000001;
  assign in_im_table_data[305] = 16'b1111000100110111;
  assign in_im_table_data[306] = 16'b1110111001011101;
  assign in_im_table_data[307] = 16'b1110110101001101;
  assign in_im_table_data[308] = 16'b1110100111110100;
  assign in_im_table_data[309] = 16'b1110100101001000;
  assign in_im_table_data[310] = 16'b1110011111010011;
  assign in_im_table_data[311] = 16'b1110011110000000;
  assign in_im_table_data[312] = 16'b1110011100001101;
  assign in_im_table_data[313] = 16'b1110011100001101;
  assign in_im_table_data[314] = 16'b1110011110000000;
  assign in_im_table_data[315] = 16'b1110011111010011;
  assign in_im_table_data[316] = 16'b1110100101001000;
  assign in_im_table_data[317] = 16'b1110100111110100;
  assign in_im_table_data[318] = 16'b1110110101001101;
  assign in_im_table_data[319] = 16'b1110111001011101;
  assign in_im_table_data[320] = 16'b1111000100110111;
  assign in_im_table_data[321] = 16'b1111001011000001;
  assign in_im_table_data[322] = 16'b1111011011011000;
  assign in_im_table_data[323] = 16'b1111100100010010;
  assign in_im_table_data[324] = 16'b1111110000101001;
  assign in_im_table_data[325] = 16'b0000000000000000;
  assign in_im_table_data[326] = 16'b0000001111010110;
  assign in_im_table_data[327] = 16'b0000011011101101;
  assign in_im_table_data[328] = 16'b0000100100100111;
  assign in_im_table_data[329] = 16'b0000110100111110;
  assign in_im_table_data[330] = 16'b0000111011001000;
  assign in_im_table_data[331] = 16'b0001000110100010;
  assign in_im_table_data[332] = 16'b0001001010110010;
  assign in_im_table_data[333] = 16'b0001011000001011;
  assign in_im_table_data[334] = 16'b0001011010110111;
  assign in_im_table_data[335] = 16'b0001100000101100;
  assign in_im_table_data[336] = 16'b0001100001111111;
  assign in_im_table_data[337] = 16'b0001100011110010;
  assign in_im_table_data[338] = 16'b0001100011110010;
  assign in_im_table_data[339] = 16'b0001100001111111;
  assign in_im_table_data[340] = 16'b0001100000101100;
  assign in_im_table_data[341] = 16'b0001011010110111;
  assign in_im_table_data[342] = 16'b0001011000001011;
  assign in_im_table_data[343] = 16'b0001001010110010;
  assign in_im_table_data[344] = 16'b0001000110100010;
  assign in_im_table_data[345] = 16'b0000111011001000;
  assign in_im_table_data[346] = 16'b0000110100111110;
  assign in_im_table_data[347] = 16'b0000100100100111;
  assign in_im_table_data[348] = 16'b0000011011101101;
  assign in_im_table_data[349] = 16'b0000001111010110;
  assign in_im_table_data[350] = 16'b0000000000000000;
  assign in_im_table_data[351] = 16'b1111110000101001;
  assign in_im_table_data[352] = 16'b1111100100010010;
  assign in_im_table_data[353] = 16'b1111011011011000;
  assign in_im_table_data[354] = 16'b1111001011000001;
  assign in_im_table_data[355] = 16'b1111000100110111;
  assign in_im_table_data[356] = 16'b1110111001011101;
  assign in_im_table_data[357] = 16'b1110110101001101;
  assign in_im_table_data[358] = 16'b1110100111110100;
  assign in_im_table_data[359] = 16'b1110100101001000;
  assign in_im_table_data[360] = 16'b1110011111010011;
  assign in_im_table_data[361] = 16'b1110011110000000;
  assign in_im_table_data[362] = 16'b1110011100001101;
  assign in_im_table_data[363] = 16'b1110011100001101;
  assign in_im_table_data[364] = 16'b1110011110000000;
  assign in_im_table_data[365] = 16'b1110011111010011;
  assign in_im_table_data[366] = 16'b1110100101001000;
  assign in_im_table_data[367] = 16'b1110100111110100;
  assign in_im_table_data[368] = 16'b1110110101001101;
  assign in_im_table_data[369] = 16'b1110111001011101;
  assign in_im_table_data[370] = 16'b1111000100110111;
  assign in_im_table_data[371] = 16'b1111001011000001;
  assign in_im_table_data[372] = 16'b1111011011011000;
  assign in_im_table_data[373] = 16'b1111100100010010;
  assign in_im_table_data[374] = 16'b1111110000101001;
  assign in_im_table_data[375] = 16'b0000000000000000;
  assign in_im_table_data[376] = 16'b0000001111010110;
  assign in_im_table_data[377] = 16'b0000011011101101;
  assign in_im_table_data[378] = 16'b0000100100100111;
  assign in_im_table_data[379] = 16'b0000110100111110;
  assign in_im_table_data[380] = 16'b0000111011001000;
  assign in_im_table_data[381] = 16'b0001000110100010;
  assign in_im_table_data[382] = 16'b0001001010110010;
  assign in_im_table_data[383] = 16'b0001011000001011;
  assign in_im_table_data[384] = 16'b0001011010110111;
  assign in_im_table_data[385] = 16'b0001100000101100;
  assign in_im_table_data[386] = 16'b0001100001111111;
  assign in_im_table_data[387] = 16'b0001100011110010;
  assign in_im_table_data[388] = 16'b0001100011110010;
  assign in_im_table_data[389] = 16'b0001100001111111;
  assign in_im_table_data[390] = 16'b0001100000101100;
  assign in_im_table_data[391] = 16'b0001011010110111;
  assign in_im_table_data[392] = 16'b0001011000001011;
  assign in_im_table_data[393] = 16'b0001001010110010;
  assign in_im_table_data[394] = 16'b0001000110100010;
  assign in_im_table_data[395] = 16'b0000111011001000;
  assign in_im_table_data[396] = 16'b0000110100111110;
  assign in_im_table_data[397] = 16'b0000100100100111;
  assign in_im_table_data[398] = 16'b0000011011101101;
  assign in_im_table_data[399] = 16'b0000001111010110;
  assign in_im_table_data[400] = 16'b0000000000000000;
  assign in_im_table_data[401] = 16'b1111110000101001;
  assign in_im_table_data[402] = 16'b1111100100010010;
  assign in_im_table_data[403] = 16'b1111011011011000;
  assign in_im_table_data[404] = 16'b1111001011000001;
  assign in_im_table_data[405] = 16'b1111000100110111;
  assign in_im_table_data[406] = 16'b1110111001011101;
  assign in_im_table_data[407] = 16'b1110110101001101;
  assign in_im_table_data[408] = 16'b1110100111110100;
  assign in_im_table_data[409] = 16'b1110100101001000;
  assign in_im_table_data[410] = 16'b1110011111010011;
  assign in_im_table_data[411] = 16'b1110011110000000;
  assign in_im_table_data[412] = 16'b1110011100001101;
  assign in_im_table_data[413] = 16'b1110011100001101;
  assign in_im_table_data[414] = 16'b1110011110000000;
  assign in_im_table_data[415] = 16'b1110011111010011;
  assign in_im_table_data[416] = 16'b1110100101001000;
  assign in_im_table_data[417] = 16'b1110100111110100;
  assign in_im_table_data[418] = 16'b1110110101001101;
  assign in_im_table_data[419] = 16'b1110111001011101;
  assign in_im_table_data[420] = 16'b1111000100110111;
  assign in_im_table_data[421] = 16'b1111001011000001;
  assign in_im_table_data[422] = 16'b1111011011011000;
  assign in_im_table_data[423] = 16'b1111100100010010;
  assign in_im_table_data[424] = 16'b1111110000101001;
  assign in_im_table_data[425] = 16'b0000000000000000;
  assign in_im_table_data[426] = 16'b0000001111010110;
  assign in_im_table_data[427] = 16'b0000011011101101;
  assign in_im_table_data[428] = 16'b0000100100100111;
  assign in_im_table_data[429] = 16'b0000110100111110;
  assign in_im_table_data[430] = 16'b0000111011001000;
  assign in_im_table_data[431] = 16'b0001000110100010;
  assign in_im_table_data[432] = 16'b0001001010110010;
  assign in_im_table_data[433] = 16'b0001011000001011;
  assign in_im_table_data[434] = 16'b0001011010110111;
  assign in_im_table_data[435] = 16'b0001100000101100;
  assign in_im_table_data[436] = 16'b0001100001111111;
  assign in_im_table_data[437] = 16'b0001100011110010;
  assign in_im_table_data[438] = 16'b0001100011110010;
  assign in_im_table_data[439] = 16'b0001100001111111;
  assign in_im_table_data[440] = 16'b0001100000101100;
  assign in_im_table_data[441] = 16'b0001011010110111;
  assign in_im_table_data[442] = 16'b0001011000001011;
  assign in_im_table_data[443] = 16'b0001001010110010;
  assign in_im_table_data[444] = 16'b0001000110100010;
  assign in_im_table_data[445] = 16'b0000111011001000;
  assign in_im_table_data[446] = 16'b0000110100111110;
  assign in_im_table_data[447] = 16'b0000100100100111;
  assign in_im_table_data[448] = 16'b0000011011101101;
  assign in_im_table_data[449] = 16'b0000001111010110;
  assign in_im_table_data[450] = 16'b0000000000000000;
  assign in_im_table_data[451] = 16'b1111110000101001;
  assign in_im_table_data[452] = 16'b1111100100010010;
  assign in_im_table_data[453] = 16'b1111011011011000;
  assign in_im_table_data[454] = 16'b1111001011000001;
  assign in_im_table_data[455] = 16'b1111000100110111;
  assign in_im_table_data[456] = 16'b1110111001011101;
  assign in_im_table_data[457] = 16'b1110110101001101;
  assign in_im_table_data[458] = 16'b1110100111110100;
  assign in_im_table_data[459] = 16'b1110100101001000;
  assign in_im_table_data[460] = 16'b1110011111010011;
  assign in_im_table_data[461] = 16'b1110011110000000;
  assign in_im_table_data[462] = 16'b1110011100001101;
  assign in_im_table_data[463] = 16'b1110011100001101;
  assign in_im_table_data[464] = 16'b1110011110000000;
  assign in_im_table_data[465] = 16'b1110011111010011;
  assign in_im_table_data[466] = 16'b1110100101001000;
  assign in_im_table_data[467] = 16'b1110100111110100;
  assign in_im_table_data[468] = 16'b1110110101001101;
  assign in_im_table_data[469] = 16'b1110111001011101;
  assign in_im_table_data[470] = 16'b1111000100110111;
  assign in_im_table_data[471] = 16'b1111001011000001;
  assign in_im_table_data[472] = 16'b1111011011011000;
  assign in_im_table_data[473] = 16'b1111100100010010;
  assign in_im_table_data[474] = 16'b1111110000101001;
  assign in_im_table_data[475] = 16'b0000000000000000;
  assign in_im_table_data[476] = 16'b0000001111010110;
  assign in_im_table_data[477] = 16'b0000011011101101;
  assign in_im_table_data[478] = 16'b0000100100100111;
  assign in_im_table_data[479] = 16'b0000110100111110;
  assign in_im_table_data[480] = 16'b0000111011001000;
  assign in_im_table_data[481] = 16'b0001000110100010;
  assign in_im_table_data[482] = 16'b0001001010110010;
  assign in_im_table_data[483] = 16'b0001011000001011;
  assign in_im_table_data[484] = 16'b0001011010110111;
  assign in_im_table_data[485] = 16'b0001100000101100;
  assign in_im_table_data[486] = 16'b0001100001111111;
  assign in_im_table_data[487] = 16'b0001100011110010;
  assign in_im_table_data[488] = 16'b0001100011110010;
  assign in_im_table_data[489] = 16'b0001100001111111;
  assign in_im_table_data[490] = 16'b0001100000101100;
  assign in_im_table_data[491] = 16'b0001011010110111;
  assign in_im_table_data[492] = 16'b0001011000001011;
  assign in_im_table_data[493] = 16'b0001001010110010;
  assign in_im_table_data[494] = 16'b0001000110100010;
  assign in_im_table_data[495] = 16'b0000111011001000;
  assign in_im_table_data[496] = 16'b0000110100111110;
  assign in_im_table_data[497] = 16'b0000100100100111;
  assign in_im_table_data[498] = 16'b0000011011101101;
  assign in_im_table_data[499] = 16'b0000001111010110;
  assign in_im_table_data[500] = 16'b1110000011111101;
  assign in_im_table_data[501] = 16'b1110001100001000;
  assign in_im_table_data[502] = 16'b1110011011001110;
  assign in_im_table_data[503] = 16'b1110101010111011;
  assign in_im_table_data[504] = 16'b1110110111001111;
  assign in_im_table_data[505] = 16'b1111000101000010;
  assign in_im_table_data[506] = 16'b1111010011000001;
  assign in_im_table_data[507] = 16'b1111100110000000;
  assign in_im_table_data[508] = 16'b1111111010100000;
  assign in_im_table_data[509] = 16'b0000001001111000;
  assign in_im_table_data[510] = 16'b0000011110100110;
  assign in_im_table_data[511] = 16'b0000110001101000;
  assign in_im_table_data[512] = 16'b0001000000100001;
  assign in_im_table_data[513] = 16'b0001001110011101;
  assign in_im_table_data[514] = 16'b0001011110111110;
  assign in_im_table_data[515] = 16'b0001101110111010;
  assign in_im_table_data[516] = 16'b0001110111110001;
  assign in_im_table_data[517] = 16'b0010000000011010;
  assign in_im_table_data[518] = 16'b0010000101010101;
  assign in_im_table_data[519] = 16'b0010001010101101;
  assign in_im_table_data[520] = 16'b0010001100011110;
  assign in_im_table_data[521] = 16'b0010010001111100;
  assign in_im_table_data[522] = 16'b0010010000110000;
  assign in_im_table_data[523] = 16'b0010001000110010;
  assign in_im_table_data[524] = 16'b0010000100011101;
  assign in_im_table_data[525] = 16'b0001111100000010;
  assign in_im_table_data[526] = 16'b0001110011110111;
  assign in_im_table_data[527] = 16'b0001100100110001;
  assign in_im_table_data[528] = 16'b0001010101000100;
  assign in_im_table_data[529] = 16'b0001001000110000;
  assign in_im_table_data[530] = 16'b0000111010111101;
  assign in_im_table_data[531] = 16'b0000101100111110;
  assign in_im_table_data[532] = 16'b0000011001111111;
  assign in_im_table_data[533] = 16'b0000000101011111;
  assign in_im_table_data[534] = 16'b1111110110000111;
  assign in_im_table_data[535] = 16'b1111100001011001;
  assign in_im_table_data[536] = 16'b1111001110010111;
  assign in_im_table_data[537] = 16'b1110111111011110;
  assign in_im_table_data[538] = 16'b1110110001100010;
  assign in_im_table_data[539] = 16'b1110100001000001;
  assign in_im_table_data[540] = 16'b1110010001000101;
  assign in_im_table_data[541] = 16'b1110001000001110;
  assign in_im_table_data[542] = 16'b1101111111100101;
  assign in_im_table_data[543] = 16'b1101111010101010;
  assign in_im_table_data[544] = 16'b1101110101010010;
  assign in_im_table_data[545] = 16'b1101110011100001;
  assign in_im_table_data[546] = 16'b1101101110000011;
  assign in_im_table_data[547] = 16'b1101101111001111;
  assign in_im_table_data[548] = 16'b1101110111001101;
  assign in_im_table_data[549] = 16'b1101111011100010;
  assign in_im_table_data[550] = 16'b1110000011111101;
  assign in_im_table_data[551] = 16'b1110001100001000;
  assign in_im_table_data[552] = 16'b1110011011001110;
  assign in_im_table_data[553] = 16'b1110101010111011;
  assign in_im_table_data[554] = 16'b1110110111001111;
  assign in_im_table_data[555] = 16'b1111000101000010;
  assign in_im_table_data[556] = 16'b1111010011000001;
  assign in_im_table_data[557] = 16'b1111100110000000;
  assign in_im_table_data[558] = 16'b1111111010100000;
  assign in_im_table_data[559] = 16'b0000001001111000;
  assign in_im_table_data[560] = 16'b0000011110100110;
  assign in_im_table_data[561] = 16'b0000110001101000;
  assign in_im_table_data[562] = 16'b0001000000100001;
  assign in_im_table_data[563] = 16'b0001001110011101;
  assign in_im_table_data[564] = 16'b0001011110111110;
  assign in_im_table_data[565] = 16'b0001101110111010;
  assign in_im_table_data[566] = 16'b0001110111110001;
  assign in_im_table_data[567] = 16'b0010000000011010;
  assign in_im_table_data[568] = 16'b0010000101010101;
  assign in_im_table_data[569] = 16'b0010001010101101;
  assign in_im_table_data[570] = 16'b0010001100011110;
  assign in_im_table_data[571] = 16'b0010010001111100;
  assign in_im_table_data[572] = 16'b0010010000110000;
  assign in_im_table_data[573] = 16'b0010001000110010;
  assign in_im_table_data[574] = 16'b0010000100011101;
  assign in_im_table_data[575] = 16'b0001111100000010;
  assign in_im_table_data[576] = 16'b0001110011110111;
  assign in_im_table_data[577] = 16'b0001100100110001;
  assign in_im_table_data[578] = 16'b0001010101000100;
  assign in_im_table_data[579] = 16'b0001001000110000;
  assign in_im_table_data[580] = 16'b0000111010111101;
  assign in_im_table_data[581] = 16'b0000101100111110;
  assign in_im_table_data[582] = 16'b0000011001111111;
  assign in_im_table_data[583] = 16'b0000000101011111;
  assign in_im_table_data[584] = 16'b1111110110000111;
  assign in_im_table_data[585] = 16'b1111100001011001;
  assign in_im_table_data[586] = 16'b1111001110010111;
  assign in_im_table_data[587] = 16'b1110111111011110;
  assign in_im_table_data[588] = 16'b1110110001100010;
  assign in_im_table_data[589] = 16'b1110100001000001;
  assign in_im_table_data[590] = 16'b1110010001000101;
  assign in_im_table_data[591] = 16'b1110001000001110;
  assign in_im_table_data[592] = 16'b1101111111100101;
  assign in_im_table_data[593] = 16'b1101111010101010;
  assign in_im_table_data[594] = 16'b1101110101010010;
  assign in_im_table_data[595] = 16'b1101110011100001;
  assign in_im_table_data[596] = 16'b1101101110000011;
  assign in_im_table_data[597] = 16'b1101101111001111;
  assign in_im_table_data[598] = 16'b1101110111001101;
  assign in_im_table_data[599] = 16'b1101111011100010;
  assign in_im_table_data[600] = 16'b1110000011111101;
  assign in_im_table_data[601] = 16'b1110001100001000;
  assign in_im_table_data[602] = 16'b1110011011001110;
  assign in_im_table_data[603] = 16'b1110101010111011;
  assign in_im_table_data[604] = 16'b1110110111001111;
  assign in_im_table_data[605] = 16'b1111000101000010;
  assign in_im_table_data[606] = 16'b1111010011000001;
  assign in_im_table_data[607] = 16'b1111100110000000;
  assign in_im_table_data[608] = 16'b1111111010100000;
  assign in_im_table_data[609] = 16'b0000001001111000;
  assign in_im_table_data[610] = 16'b0000011110100110;
  assign in_im_table_data[611] = 16'b0000110001101000;
  assign in_im_table_data[612] = 16'b0001000000100001;
  assign in_im_table_data[613] = 16'b0001001110011101;
  assign in_im_table_data[614] = 16'b0001011110111110;
  assign in_im_table_data[615] = 16'b0001101110111010;
  assign in_im_table_data[616] = 16'b0001110111110001;
  assign in_im_table_data[617] = 16'b0010000000011010;
  assign in_im_table_data[618] = 16'b0010000101010101;
  assign in_im_table_data[619] = 16'b0010001010101101;
  assign in_im_table_data[620] = 16'b0010001100011110;
  assign in_im_table_data[621] = 16'b0010010001111100;
  assign in_im_table_data[622] = 16'b0010010000110000;
  assign in_im_table_data[623] = 16'b0010001000110010;
  assign in_im_table_data[624] = 16'b0010000100011101;
  assign in_im_table_data[625] = 16'b0001111100000010;
  assign in_im_table_data[626] = 16'b0001110011110111;
  assign in_im_table_data[627] = 16'b0001100100110001;
  assign in_im_table_data[628] = 16'b0001010101000100;
  assign in_im_table_data[629] = 16'b0001001000110000;
  assign in_im_table_data[630] = 16'b0000111010111101;
  assign in_im_table_data[631] = 16'b0000101100111110;
  assign in_im_table_data[632] = 16'b0000011001111111;
  assign in_im_table_data[633] = 16'b0000000101011111;
  assign in_im_table_data[634] = 16'b1111110110000111;
  assign in_im_table_data[635] = 16'b1111100001011001;
  assign in_im_table_data[636] = 16'b1111001110010111;
  assign in_im_table_data[637] = 16'b1110111111011110;
  assign in_im_table_data[638] = 16'b1110110001100010;
  assign in_im_table_data[639] = 16'b1110100001000001;
  assign in_im_table_data[640] = 16'b1110010001000101;
  assign in_im_table_data[641] = 16'b1110001000001110;
  assign in_im_table_data[642] = 16'b1101111111100101;
  assign in_im_table_data[643] = 16'b1101111010101010;
  assign in_im_table_data[644] = 16'b1101110101010010;
  assign in_im_table_data[645] = 16'b1101110011100001;
  assign in_im_table_data[646] = 16'b1101101110000011;
  assign in_im_table_data[647] = 16'b1101101111001111;
  assign in_im_table_data[648] = 16'b1101110111001101;
  assign in_im_table_data[649] = 16'b1101111011100010;
  assign in_im_table_data[650] = 16'b1110000011111101;
  assign in_im_table_data[651] = 16'b1110001100001000;
  assign in_im_table_data[652] = 16'b1110011011001110;
  assign in_im_table_data[653] = 16'b1110101010111011;
  assign in_im_table_data[654] = 16'b1110110111001111;
  assign in_im_table_data[655] = 16'b1111000101000010;
  assign in_im_table_data[656] = 16'b1111010011000001;
  assign in_im_table_data[657] = 16'b1111100110000000;
  assign in_im_table_data[658] = 16'b1111111010100000;
  assign in_im_table_data[659] = 16'b0000001001111000;
  assign in_im_table_data[660] = 16'b0000011110100110;
  assign in_im_table_data[661] = 16'b0000110001101000;
  assign in_im_table_data[662] = 16'b0001000000100001;
  assign in_im_table_data[663] = 16'b0001001110011101;
  assign in_im_table_data[664] = 16'b0001011110111110;
  assign in_im_table_data[665] = 16'b0001101110111010;
  assign in_im_table_data[666] = 16'b0001110111110001;
  assign in_im_table_data[667] = 16'b0010000000011010;
  assign in_im_table_data[668] = 16'b0010000101010101;
  assign in_im_table_data[669] = 16'b0010001010101101;
  assign in_im_table_data[670] = 16'b0010001100011110;
  assign in_im_table_data[671] = 16'b0010010001111100;
  assign in_im_table_data[672] = 16'b0010010000110000;
  assign in_im_table_data[673] = 16'b0010001000110010;
  assign in_im_table_data[674] = 16'b0010000100011101;
  assign in_im_table_data[675] = 16'b0001111100000010;
  assign in_im_table_data[676] = 16'b0001110011110111;
  assign in_im_table_data[677] = 16'b0001100100110001;
  assign in_im_table_data[678] = 16'b0001010101000100;
  assign in_im_table_data[679] = 16'b0001001000110000;
  assign in_im_table_data[680] = 16'b0000111010111101;
  assign in_im_table_data[681] = 16'b0000101100111110;
  assign in_im_table_data[682] = 16'b0000011001111111;
  assign in_im_table_data[683] = 16'b0000000101011111;
  assign in_im_table_data[684] = 16'b1111110110000111;
  assign in_im_table_data[685] = 16'b1111100001011001;
  assign in_im_table_data[686] = 16'b1111001110010111;
  assign in_im_table_data[687] = 16'b1110111111011110;
  assign in_im_table_data[688] = 16'b1110110001100010;
  assign in_im_table_data[689] = 16'b1110100001000001;
  assign in_im_table_data[690] = 16'b1110010001000101;
  assign in_im_table_data[691] = 16'b1110001000001110;
  assign in_im_table_data[692] = 16'b1101111111100101;
  assign in_im_table_data[693] = 16'b1101111010101010;
  assign in_im_table_data[694] = 16'b1101110101010010;
  assign in_im_table_data[695] = 16'b1101110011100001;
  assign in_im_table_data[696] = 16'b1101101110000011;
  assign in_im_table_data[697] = 16'b1101101111001111;
  assign in_im_table_data[698] = 16'b1101110111001101;
  assign in_im_table_data[699] = 16'b1101111011100010;
  assign in_im_table_data[700] = 16'b1110000011111101;
  assign in_im_table_data[701] = 16'b1110001100001000;
  assign in_im_table_data[702] = 16'b1110011011001110;
  assign in_im_table_data[703] = 16'b1110101010111011;
  assign in_im_table_data[704] = 16'b1110110111001111;
  assign in_im_table_data[705] = 16'b1111000101000010;
  assign in_im_table_data[706] = 16'b1111010011000001;
  assign in_im_table_data[707] = 16'b1111100110000000;
  assign in_im_table_data[708] = 16'b1111111010100000;
  assign in_im_table_data[709] = 16'b0000001001111000;
  assign in_im_table_data[710] = 16'b0000011110100110;
  assign in_im_table_data[711] = 16'b0000110001101000;
  assign in_im_table_data[712] = 16'b0001000000100001;
  assign in_im_table_data[713] = 16'b0001001110011101;
  assign in_im_table_data[714] = 16'b0001011110111110;
  assign in_im_table_data[715] = 16'b0001101110111010;
  assign in_im_table_data[716] = 16'b0001110111110001;
  assign in_im_table_data[717] = 16'b0010000000011010;
  assign in_im_table_data[718] = 16'b0010000101010101;
  assign in_im_table_data[719] = 16'b0010001010101101;
  assign in_im_table_data[720] = 16'b0010001100011110;
  assign in_im_table_data[721] = 16'b0010010001111100;
  assign in_im_table_data[722] = 16'b0010010000110000;
  assign in_im_table_data[723] = 16'b0010001000110010;
  assign in_im_table_data[724] = 16'b0010000100011101;
  assign in_im_table_data[725] = 16'b0001111100000010;
  assign in_im_table_data[726] = 16'b0001110011110111;
  assign in_im_table_data[727] = 16'b0001100100110001;
  assign in_im_table_data[728] = 16'b0001010101000100;
  assign in_im_table_data[729] = 16'b0001001000110000;
  assign in_im_table_data[730] = 16'b0000111010111101;
  assign in_im_table_data[731] = 16'b0000101100111110;
  assign in_im_table_data[732] = 16'b0000011001111111;
  assign in_im_table_data[733] = 16'b0000000101011111;
  assign in_im_table_data[734] = 16'b1111110110000111;
  assign in_im_table_data[735] = 16'b1111100001011001;
  assign in_im_table_data[736] = 16'b1111001110010111;
  assign in_im_table_data[737] = 16'b1110111111011110;
  assign in_im_table_data[738] = 16'b1110110001100010;
  assign in_im_table_data[739] = 16'b1110100001000001;
  assign in_im_table_data[740] = 16'b1110010001000101;
  assign in_im_table_data[741] = 16'b1110001000001110;
  assign in_im_table_data[742] = 16'b1101111111100101;
  assign in_im_table_data[743] = 16'b1101111010101010;
  assign in_im_table_data[744] = 16'b1101110101010010;
  assign in_im_table_data[745] = 16'b1101110011100001;
  assign in_im_table_data[746] = 16'b1101101110000011;
  assign in_im_table_data[747] = 16'b1101101111001111;
  assign in_im_table_data[748] = 16'b1101110111001101;
  assign in_im_table_data[749] = 16'b1101111011100010;
  assign in_im_table_data[750] = 16'b0000001010011100;
  assign in_im_table_data[751] = 16'b0000000110000000;
  assign in_im_table_data[752] = 16'b0000000111110111;
  assign in_im_table_data[753] = 16'b0000000110111100;
  assign in_im_table_data[754] = 16'b0000001001001110;
  assign in_im_table_data[755] = 16'b0000001001001100;
  assign in_im_table_data[756] = 16'b0000001110101010;
  assign in_im_table_data[757] = 16'b0000001111010001;
  assign in_im_table_data[758] = 16'b0000001010011000;
  assign in_im_table_data[759] = 16'b0000001011111010;
  assign in_im_table_data[760] = 16'b0000001010010001;
  assign in_im_table_data[761] = 16'b0000001111011001;
  assign in_im_table_data[762] = 16'b0000001110010010;
  assign in_im_table_data[763] = 16'b0000001001011100;
  assign in_im_table_data[764] = 16'b0000001000011110;
  assign in_im_table_data[765] = 16'b0000000111010111;
  assign in_im_table_data[766] = 16'b0000000110010111;
  assign in_im_table_data[767] = 16'b0000000110101001;
  assign in_im_table_data[768] = 16'b0000000101011111;
  assign in_im_table_data[769] = 16'b0000001001011110;
  assign in_im_table_data[770] = 16'b0000001000000000;
  assign in_im_table_data[771] = 16'b0000000001111100;
  assign in_im_table_data[772] = 16'b1111111111110001;
  assign in_im_table_data[773] = 16'b1111111101001010;
  assign in_im_table_data[774] = 16'b1111110111100000;
  assign in_im_table_data[775] = 16'b1111110101100011;
  assign in_im_table_data[776] = 16'b1111111001111111;
  assign in_im_table_data[777] = 16'b1111111000001000;
  assign in_im_table_data[778] = 16'b1111111001000011;
  assign in_im_table_data[779] = 16'b1111110110110001;
  assign in_im_table_data[780] = 16'b1111110110110011;
  assign in_im_table_data[781] = 16'b1111110001010101;
  assign in_im_table_data[782] = 16'b1111110000101110;
  assign in_im_table_data[783] = 16'b1111110101100111;
  assign in_im_table_data[784] = 16'b1111110100000101;
  assign in_im_table_data[785] = 16'b1111110101101110;
  assign in_im_table_data[786] = 16'b1111110000100110;
  assign in_im_table_data[787] = 16'b1111110001101101;
  assign in_im_table_data[788] = 16'b1111110110100011;
  assign in_im_table_data[789] = 16'b1111110111100001;
  assign in_im_table_data[790] = 16'b1111111000101000;
  assign in_im_table_data[791] = 16'b1111111001101000;
  assign in_im_table_data[792] = 16'b1111111001010110;
  assign in_im_table_data[793] = 16'b1111111010100000;
  assign in_im_table_data[794] = 16'b1111110110100001;
  assign in_im_table_data[795] = 16'b1111110111111111;
  assign in_im_table_data[796] = 16'b1111111110000011;
  assign in_im_table_data[797] = 16'b0000000000001110;
  assign in_im_table_data[798] = 16'b0000000010110101;
  assign in_im_table_data[799] = 16'b0000001000011111;
  assign in_im_table_data[800] = 16'b0000001010011100;
  assign in_im_table_data[801] = 16'b0000000110000000;
  assign in_im_table_data[802] = 16'b0000000111110111;
  assign in_im_table_data[803] = 16'b0000000110111100;
  assign in_im_table_data[804] = 16'b0000001001001110;
  assign in_im_table_data[805] = 16'b0000001001001100;
  assign in_im_table_data[806] = 16'b0000001110101010;
  assign in_im_table_data[807] = 16'b0000001111010001;
  assign in_im_table_data[808] = 16'b0000001010011000;
  assign in_im_table_data[809] = 16'b0000001011111010;
  assign in_im_table_data[810] = 16'b0000001010010001;
  assign in_im_table_data[811] = 16'b0000001111011001;
  assign in_im_table_data[812] = 16'b0000001110010010;
  assign in_im_table_data[813] = 16'b0000001001011100;
  assign in_im_table_data[814] = 16'b0000001000011110;
  assign in_im_table_data[815] = 16'b0000000111010111;
  assign in_im_table_data[816] = 16'b0000000110010111;
  assign in_im_table_data[817] = 16'b0000000110101001;
  assign in_im_table_data[818] = 16'b0000000101011111;
  assign in_im_table_data[819] = 16'b0000001001011110;
  assign in_im_table_data[820] = 16'b0000001000000000;
  assign in_im_table_data[821] = 16'b0000000001111100;
  assign in_im_table_data[822] = 16'b1111111111110001;
  assign in_im_table_data[823] = 16'b1111111101001010;
  assign in_im_table_data[824] = 16'b1111110111100000;
  assign in_im_table_data[825] = 16'b1111110101100011;
  assign in_im_table_data[826] = 16'b1111111001111111;
  assign in_im_table_data[827] = 16'b1111111000001000;
  assign in_im_table_data[828] = 16'b1111111001000011;
  assign in_im_table_data[829] = 16'b1111110110110001;
  assign in_im_table_data[830] = 16'b1111110110110011;
  assign in_im_table_data[831] = 16'b1111110001010101;
  assign in_im_table_data[832] = 16'b1111110000101110;
  assign in_im_table_data[833] = 16'b1111110101100111;
  assign in_im_table_data[834] = 16'b1111110100000101;
  assign in_im_table_data[835] = 16'b1111110101101110;
  assign in_im_table_data[836] = 16'b1111110000100110;
  assign in_im_table_data[837] = 16'b1111110001101101;
  assign in_im_table_data[838] = 16'b1111110110100011;
  assign in_im_table_data[839] = 16'b1111110111100001;
  assign in_im_table_data[840] = 16'b1111111000101000;
  assign in_im_table_data[841] = 16'b1111111001101000;
  assign in_im_table_data[842] = 16'b1111111001010110;
  assign in_im_table_data[843] = 16'b1111111010100000;
  assign in_im_table_data[844] = 16'b1111110110100001;
  assign in_im_table_data[845] = 16'b1111110111111111;
  assign in_im_table_data[846] = 16'b1111111110000011;
  assign in_im_table_data[847] = 16'b0000000000001110;
  assign in_im_table_data[848] = 16'b0000000010110101;
  assign in_im_table_data[849] = 16'b0000001000011111;
  assign in_im_table_data[850] = 16'b0000001010011100;
  assign in_im_table_data[851] = 16'b0000000110000000;
  assign in_im_table_data[852] = 16'b0000000111110111;
  assign in_im_table_data[853] = 16'b0000000110111100;
  assign in_im_table_data[854] = 16'b0000001001001110;
  assign in_im_table_data[855] = 16'b0000001001001100;
  assign in_im_table_data[856] = 16'b0000001110101010;
  assign in_im_table_data[857] = 16'b0000001111010001;
  assign in_im_table_data[858] = 16'b0000001010011000;
  assign in_im_table_data[859] = 16'b0000001011111010;
  assign in_im_table_data[860] = 16'b0000001010010001;
  assign in_im_table_data[861] = 16'b0000001111011001;
  assign in_im_table_data[862] = 16'b0000001110010010;
  assign in_im_table_data[863] = 16'b0000001001011100;
  assign in_im_table_data[864] = 16'b0000001000011110;
  assign in_im_table_data[865] = 16'b0000000111010111;
  assign in_im_table_data[866] = 16'b0000000110010111;
  assign in_im_table_data[867] = 16'b0000000110101001;
  assign in_im_table_data[868] = 16'b0000000101011111;
  assign in_im_table_data[869] = 16'b0000001001011110;
  assign in_im_table_data[870] = 16'b0000001000000000;
  assign in_im_table_data[871] = 16'b0000000001111100;
  assign in_im_table_data[872] = 16'b1111111111110001;
  assign in_im_table_data[873] = 16'b1111111101001010;
  assign in_im_table_data[874] = 16'b1111110111100000;
  assign in_im_table_data[875] = 16'b1111110101100011;
  assign in_im_table_data[876] = 16'b1111111001111111;
  assign in_im_table_data[877] = 16'b1111111000001000;
  assign in_im_table_data[878] = 16'b1111111001000011;
  assign in_im_table_data[879] = 16'b1111110110110001;
  assign in_im_table_data[880] = 16'b1111110110110011;
  assign in_im_table_data[881] = 16'b1111110001010101;
  assign in_im_table_data[882] = 16'b1111110000101110;
  assign in_im_table_data[883] = 16'b1111110101100111;
  assign in_im_table_data[884] = 16'b1111110100000101;
  assign in_im_table_data[885] = 16'b1111110101101110;
  assign in_im_table_data[886] = 16'b1111110000100110;
  assign in_im_table_data[887] = 16'b1111110001101101;
  assign in_im_table_data[888] = 16'b1111110110100011;
  assign in_im_table_data[889] = 16'b1111110111100001;
  assign in_im_table_data[890] = 16'b1111111000101000;
  assign in_im_table_data[891] = 16'b1111111001101000;
  assign in_im_table_data[892] = 16'b1111111001010110;
  assign in_im_table_data[893] = 16'b1111111010100000;
  assign in_im_table_data[894] = 16'b1111110110100001;
  assign in_im_table_data[895] = 16'b1111110111111111;
  assign in_im_table_data[896] = 16'b1111111110000011;
  assign in_im_table_data[897] = 16'b0000000000001110;
  assign in_im_table_data[898] = 16'b0000000010110101;
  assign in_im_table_data[899] = 16'b0000001000011111;
  assign in_im_table_data[900] = 16'b0000001010011100;
  assign in_im_table_data[901] = 16'b0000000110000000;
  assign in_im_table_data[902] = 16'b0000000111110111;
  assign in_im_table_data[903] = 16'b0000000110111100;
  assign in_im_table_data[904] = 16'b0000001001001110;
  assign in_im_table_data[905] = 16'b0000001001001100;
  assign in_im_table_data[906] = 16'b0000001110101010;
  assign in_im_table_data[907] = 16'b0000001111010001;
  assign in_im_table_data[908] = 16'b0000001010011000;
  assign in_im_table_data[909] = 16'b0000001011111010;
  assign in_im_table_data[910] = 16'b0000001010010001;
  assign in_im_table_data[911] = 16'b0000001111011001;
  assign in_im_table_data[912] = 16'b0000001110010010;
  assign in_im_table_data[913] = 16'b0000001001011100;
  assign in_im_table_data[914] = 16'b0000001000011110;
  assign in_im_table_data[915] = 16'b0000000111010111;
  assign in_im_table_data[916] = 16'b0000000110010111;
  assign in_im_table_data[917] = 16'b0000000110101001;
  assign in_im_table_data[918] = 16'b0000000101011111;
  assign in_im_table_data[919] = 16'b0000001001011110;
  assign in_im_table_data[920] = 16'b0000001000000000;
  assign in_im_table_data[921] = 16'b0000000001111100;
  assign in_im_table_data[922] = 16'b1111111111110001;
  assign in_im_table_data[923] = 16'b1111111101001010;
  assign in_im_table_data[924] = 16'b1111110111100000;
  assign in_im_table_data[925] = 16'b1111110101100011;
  assign in_im_table_data[926] = 16'b1111111001111111;
  assign in_im_table_data[927] = 16'b1111111000001000;
  assign in_im_table_data[928] = 16'b1111111001000011;
  assign in_im_table_data[929] = 16'b1111110110110001;
  assign in_im_table_data[930] = 16'b1111110110110011;
  assign in_im_table_data[931] = 16'b1111110001010101;
  assign in_im_table_data[932] = 16'b1111110000101110;
  assign in_im_table_data[933] = 16'b1111110101100111;
  assign in_im_table_data[934] = 16'b1111110100000101;
  assign in_im_table_data[935] = 16'b1111110101101110;
  assign in_im_table_data[936] = 16'b1111110000100110;
  assign in_im_table_data[937] = 16'b1111110001101101;
  assign in_im_table_data[938] = 16'b1111110110100011;
  assign in_im_table_data[939] = 16'b1111110111100001;
  assign in_im_table_data[940] = 16'b1111111000101000;
  assign in_im_table_data[941] = 16'b1111111001101000;
  assign in_im_table_data[942] = 16'b1111111001010110;
  assign in_im_table_data[943] = 16'b1111111010100000;
  assign in_im_table_data[944] = 16'b1111110110100001;
  assign in_im_table_data[945] = 16'b1111110111111111;
  assign in_im_table_data[946] = 16'b1111111110000011;
  assign in_im_table_data[947] = 16'b0000000000001110;
  assign in_im_table_data[948] = 16'b0000000010110101;
  assign in_im_table_data[949] = 16'b0000001000011111;
  assign in_im_table_data[950] = 16'b0000001010011100;
  assign in_im_table_data[951] = 16'b0000000110000000;
  assign in_im_table_data[952] = 16'b0000000111110111;
  assign in_im_table_data[953] = 16'b0000000110111100;
  assign in_im_table_data[954] = 16'b0000001001001110;
  assign in_im_table_data[955] = 16'b0000001001001100;
  assign in_im_table_data[956] = 16'b0000001110101010;
  assign in_im_table_data[957] = 16'b0000001111010001;
  assign in_im_table_data[958] = 16'b0000001010011000;
  assign in_im_table_data[959] = 16'b0000001011111010;
  assign in_im_table_data[960] = 16'b0000001010010001;
  assign in_im_table_data[961] = 16'b0000001111011001;
  assign in_im_table_data[962] = 16'b0000001110010010;
  assign in_im_table_data[963] = 16'b0000001001011100;
  assign in_im_table_data[964] = 16'b0000001000011110;
  assign in_im_table_data[965] = 16'b0000000111010111;
  assign in_im_table_data[966] = 16'b0000000110010111;
  assign in_im_table_data[967] = 16'b0000000110101001;
  assign in_im_table_data[968] = 16'b0000000101011111;
  assign in_im_table_data[969] = 16'b0000001001011110;
  assign in_im_table_data[970] = 16'b0000001000000000;
  assign in_im_table_data[971] = 16'b0000000001111100;
  assign in_im_table_data[972] = 16'b1111111111110001;
  assign in_im_table_data[973] = 16'b1111111101001010;
  assign in_im_table_data[974] = 16'b1111110111100000;
  assign in_im_table_data[975] = 16'b1111110101100011;
  assign in_im_table_data[976] = 16'b1111111001111111;
  assign in_im_table_data[977] = 16'b1111111000001000;
  assign in_im_table_data[978] = 16'b1111111001000011;
  assign in_im_table_data[979] = 16'b1111110110110001;
  assign in_im_table_data[980] = 16'b1111110110110011;
  assign in_im_table_data[981] = 16'b1111110001010101;
  assign in_im_table_data[982] = 16'b1111110000101110;
  assign in_im_table_data[983] = 16'b1111110101100111;
  assign in_im_table_data[984] = 16'b1111110100000101;
  assign in_im_table_data[985] = 16'b1111110101101110;
  assign in_im_table_data[986] = 16'b1111110000100110;
  assign in_im_table_data[987] = 16'b1111110001101101;
  assign in_im_table_data[988] = 16'b1111110110100011;
  assign in_im_table_data[989] = 16'b1111110111100001;
  assign in_im_table_data[990] = 16'b1111111000101000;
  assign in_im_table_data[991] = 16'b1111111001101000;
  assign in_im_table_data[992] = 16'b1111111001010110;
  assign in_im_table_data[993] = 16'b1111111010100000;
  assign in_im_table_data[994] = 16'b1111110110100001;
  assign in_im_table_data[995] = 16'b1111110111111111;
  assign in_im_table_data[996] = 16'b1111111110000011;
  assign in_im_table_data[997] = 16'b0000000000001110;
  assign in_im_table_data[998] = 16'b0000000010110101;
  assign in_im_table_data[999] = 16'b0000001000011111;
  assign in_im_table_data[1000] = 16'b1111110111100000;
  assign in_im_1 = in_im_table_data[Data_Type_Conversion1_out1_addr];



  assign rawData_in_im = in_im_1;



  // holdData reg for Data_Type_Conversion1_out1
  always @(posedge clk)
    begin : stimuli_Data_Type_Conversion1_out1
      if (reset_x) begin
        holdData_in_im <= 16'bx;
      end
      else begin
        holdData_in_im <= rawData_in_im;
      end
    end

  always @(rawData_in_im or rdEnb)
    begin : stimuli_Data_Type_Conversion1_out1_1
      if (rdEnb == 1'b0) begin
        in_im_offset <= holdData_in_im;
      end
      else begin
        in_im_offset <= rawData_in_im;
      end
    end

  assign #2 in_im_2 = in_im_offset;

  assign Data_Type_Conversion1_out1_active = Data_Type_Conversion1_out1_addr != 10'b1111101000;



  assign Data_Type_Conversion1_out1_enb = Data_Type_Conversion1_out1_active & (rdEnb & tb_enb_delay);



  // Count limited, Unsigned Counter
  //  initial value   = 0
  //  step value      = 1
  //  count to value  = 1000
  always @(posedge clk)
    begin : DataTypeConversion1_process
      if (reset_x == 1'b1) begin
        Data_Type_Conversion1_out1_addr <= 10'b0000000000;
      end
      else begin
        if (Data_Type_Conversion1_out1_enb) begin
          if (Data_Type_Conversion1_out1_addr >= 10'b1111101000) begin
            Data_Type_Conversion1_out1_addr <= 10'b0000000000;
          end
          else begin
            Data_Type_Conversion1_out1_addr <= Data_Type_Conversion1_out1_addr + 10'b0000000001;
          end
        end
      end
    end



  // Data source for in_re
  assign in_re_table_data[0] = 16'b0100111111111111;
  assign in_re_table_data[1] = 16'b0101000000000000;
  assign in_re_table_data[2] = 16'b0100110111111111;
  assign in_re_table_data[3] = 16'b0100100111111111;
  assign in_re_table_data[4] = 16'b0100010111111111;
  assign in_re_table_data[5] = 16'b0100000000000000;
  assign in_re_table_data[6] = 16'b0011100111111111;
  assign in_re_table_data[7] = 16'b0011000111111111;
  assign in_re_table_data[8] = 16'b0010100111111111;
  assign in_re_table_data[9] = 16'b0010001000000000;
  assign in_re_table_data[10] = 16'b0001011111111111;
  assign in_re_table_data[11] = 16'b0000111000000000;
  assign in_re_table_data[12] = 16'b0000011000000000;
  assign in_re_table_data[13] = 16'b1111101000000000;
  assign in_re_table_data[14] = 16'b1111001000000000;
  assign in_re_table_data[15] = 16'b1110100000000000;
  assign in_re_table_data[16] = 16'b1101111000000000;
  assign in_re_table_data[17] = 16'b1101011000000000;
  assign in_re_table_data[18] = 16'b1100111000000000;
  assign in_re_table_data[19] = 16'b1100011000000000;
  assign in_re_table_data[20] = 16'b1100000000000000;
  assign in_re_table_data[21] = 16'b1011101000000000;
  assign in_re_table_data[22] = 16'b1011011000000000;
  assign in_re_table_data[23] = 16'b1011001000000000;
  assign in_re_table_data[24] = 16'b1011000000000000;
  assign in_re_table_data[25] = 16'b1011000000000000;
  assign in_re_table_data[26] = 16'b1011000000000000;
  assign in_re_table_data[27] = 16'b1011001000000000;
  assign in_re_table_data[28] = 16'b1011011000000000;
  assign in_re_table_data[29] = 16'b1011101000000000;
  assign in_re_table_data[30] = 16'b1100000000000000;
  assign in_re_table_data[31] = 16'b1100011000000000;
  assign in_re_table_data[32] = 16'b1100111000000000;
  assign in_re_table_data[33] = 16'b1101010111111111;
  assign in_re_table_data[34] = 16'b1101111000000000;
  assign in_re_table_data[35] = 16'b1110011111111111;
  assign in_re_table_data[36] = 16'b1111000111111111;
  assign in_re_table_data[37] = 16'b1111101000000000;
  assign in_re_table_data[38] = 16'b0000010111111111;
  assign in_re_table_data[39] = 16'b0000110111111111;
  assign in_re_table_data[40] = 16'b0001011111111111;
  assign in_re_table_data[41] = 16'b0010000111111111;
  assign in_re_table_data[42] = 16'b0010101000000000;
  assign in_re_table_data[43] = 16'b0011000111111111;
  assign in_re_table_data[44] = 16'b0011101000000000;
  assign in_re_table_data[45] = 16'b0100000000000000;
  assign in_re_table_data[46] = 16'b0100011000000000;
  assign in_re_table_data[47] = 16'b0100100111111111;
  assign in_re_table_data[48] = 16'b0100111000000000;
  assign in_re_table_data[49] = 16'b0101000000000000;
  assign in_re_table_data[50] = 16'b0100111111111111;
  assign in_re_table_data[51] = 16'b0101000000000000;
  assign in_re_table_data[52] = 16'b0100110111111111;
  assign in_re_table_data[53] = 16'b0100100111111111;
  assign in_re_table_data[54] = 16'b0100010111111111;
  assign in_re_table_data[55] = 16'b0100000000000000;
  assign in_re_table_data[56] = 16'b0011100111111111;
  assign in_re_table_data[57] = 16'b0011000111111111;
  assign in_re_table_data[58] = 16'b0010100111111111;
  assign in_re_table_data[59] = 16'b0010001000000000;
  assign in_re_table_data[60] = 16'b0001011111111111;
  assign in_re_table_data[61] = 16'b0000111000000000;
  assign in_re_table_data[62] = 16'b0000011000000000;
  assign in_re_table_data[63] = 16'b1111101000000000;
  assign in_re_table_data[64] = 16'b1111001000000000;
  assign in_re_table_data[65] = 16'b1110100000000000;
  assign in_re_table_data[66] = 16'b1101111000000000;
  assign in_re_table_data[67] = 16'b1101011000000000;
  assign in_re_table_data[68] = 16'b1100111000000000;
  assign in_re_table_data[69] = 16'b1100011000000000;
  assign in_re_table_data[70] = 16'b1100000000000000;
  assign in_re_table_data[71] = 16'b1011101000000000;
  assign in_re_table_data[72] = 16'b1011011000000000;
  assign in_re_table_data[73] = 16'b1011001000000000;
  assign in_re_table_data[74] = 16'b1011000000000000;
  assign in_re_table_data[75] = 16'b1011000000000000;
  assign in_re_table_data[76] = 16'b1011000000000000;
  assign in_re_table_data[77] = 16'b1011001000000000;
  assign in_re_table_data[78] = 16'b1011011000000000;
  assign in_re_table_data[79] = 16'b1011101000000000;
  assign in_re_table_data[80] = 16'b1100000000000000;
  assign in_re_table_data[81] = 16'b1100011000000000;
  assign in_re_table_data[82] = 16'b1100111000000000;
  assign in_re_table_data[83] = 16'b1101010111111111;
  assign in_re_table_data[84] = 16'b1101111000000000;
  assign in_re_table_data[85] = 16'b1110011111111111;
  assign in_re_table_data[86] = 16'b1111000111111111;
  assign in_re_table_data[87] = 16'b1111101000000000;
  assign in_re_table_data[88] = 16'b0000010111111111;
  assign in_re_table_data[89] = 16'b0000110111111111;
  assign in_re_table_data[90] = 16'b0001011111111111;
  assign in_re_table_data[91] = 16'b0010000111111111;
  assign in_re_table_data[92] = 16'b0010101000000000;
  assign in_re_table_data[93] = 16'b0011000111111111;
  assign in_re_table_data[94] = 16'b0011101000000000;
  assign in_re_table_data[95] = 16'b0100000000000000;
  assign in_re_table_data[96] = 16'b0100011000000000;
  assign in_re_table_data[97] = 16'b0100100111111111;
  assign in_re_table_data[98] = 16'b0100111000000000;
  assign in_re_table_data[99] = 16'b0101000000000000;
  assign in_re_table_data[100] = 16'b0100111111111111;
  assign in_re_table_data[101] = 16'b0101000000000000;
  assign in_re_table_data[102] = 16'b0100110111111111;
  assign in_re_table_data[103] = 16'b0100100111111111;
  assign in_re_table_data[104] = 16'b0100010111111111;
  assign in_re_table_data[105] = 16'b0100000000000000;
  assign in_re_table_data[106] = 16'b0011100111111111;
  assign in_re_table_data[107] = 16'b0011000111111111;
  assign in_re_table_data[108] = 16'b0010100111111111;
  assign in_re_table_data[109] = 16'b0010001000000000;
  assign in_re_table_data[110] = 16'b0001011111111111;
  assign in_re_table_data[111] = 16'b0000111000000000;
  assign in_re_table_data[112] = 16'b0000011000000000;
  assign in_re_table_data[113] = 16'b1111101000000000;
  assign in_re_table_data[114] = 16'b1111001000000000;
  assign in_re_table_data[115] = 16'b1110100000000000;
  assign in_re_table_data[116] = 16'b1101111000000000;
  assign in_re_table_data[117] = 16'b1101011000000000;
  assign in_re_table_data[118] = 16'b1100111000000000;
  assign in_re_table_data[119] = 16'b1100011000000000;
  assign in_re_table_data[120] = 16'b1100000000000000;
  assign in_re_table_data[121] = 16'b1011101000000000;
  assign in_re_table_data[122] = 16'b1011011000000000;
  assign in_re_table_data[123] = 16'b1011001000000000;
  assign in_re_table_data[124] = 16'b1011000000000000;
  assign in_re_table_data[125] = 16'b1011000000000000;
  assign in_re_table_data[126] = 16'b1011000000000000;
  assign in_re_table_data[127] = 16'b1011001000000000;
  assign in_re_table_data[128] = 16'b1011011000000000;
  assign in_re_table_data[129] = 16'b1011101000000000;
  assign in_re_table_data[130] = 16'b1100000000000000;
  assign in_re_table_data[131] = 16'b1100011000000000;
  assign in_re_table_data[132] = 16'b1100111000000000;
  assign in_re_table_data[133] = 16'b1101010111111111;
  assign in_re_table_data[134] = 16'b1101111000000000;
  assign in_re_table_data[135] = 16'b1110011111111111;
  assign in_re_table_data[136] = 16'b1111000111111111;
  assign in_re_table_data[137] = 16'b1111101000000000;
  assign in_re_table_data[138] = 16'b0000010111111111;
  assign in_re_table_data[139] = 16'b0000110111111111;
  assign in_re_table_data[140] = 16'b0001011111111111;
  assign in_re_table_data[141] = 16'b0010000111111111;
  assign in_re_table_data[142] = 16'b0010101000000000;
  assign in_re_table_data[143] = 16'b0011000111111111;
  assign in_re_table_data[144] = 16'b0011101000000000;
  assign in_re_table_data[145] = 16'b0100000000000000;
  assign in_re_table_data[146] = 16'b0100011000000000;
  assign in_re_table_data[147] = 16'b0100100111111111;
  assign in_re_table_data[148] = 16'b0100111000000000;
  assign in_re_table_data[149] = 16'b0101000000000000;
  assign in_re_table_data[150] = 16'b0100111111111111;
  assign in_re_table_data[151] = 16'b0101000000000000;
  assign in_re_table_data[152] = 16'b0100110111111111;
  assign in_re_table_data[153] = 16'b0100100111111111;
  assign in_re_table_data[154] = 16'b0100010111111111;
  assign in_re_table_data[155] = 16'b0100000000000000;
  assign in_re_table_data[156] = 16'b0011100111111111;
  assign in_re_table_data[157] = 16'b0011000111111111;
  assign in_re_table_data[158] = 16'b0010100111111111;
  assign in_re_table_data[159] = 16'b0010001000000000;
  assign in_re_table_data[160] = 16'b0001011111111111;
  assign in_re_table_data[161] = 16'b0000111000000000;
  assign in_re_table_data[162] = 16'b0000011000000000;
  assign in_re_table_data[163] = 16'b1111101000000000;
  assign in_re_table_data[164] = 16'b1111001000000000;
  assign in_re_table_data[165] = 16'b1110100000000000;
  assign in_re_table_data[166] = 16'b1101111000000000;
  assign in_re_table_data[167] = 16'b1101011000000000;
  assign in_re_table_data[168] = 16'b1100111000000000;
  assign in_re_table_data[169] = 16'b1100011000000000;
  assign in_re_table_data[170] = 16'b1100000000000000;
  assign in_re_table_data[171] = 16'b1011101000000000;
  assign in_re_table_data[172] = 16'b1011011000000000;
  assign in_re_table_data[173] = 16'b1011001000000000;
  assign in_re_table_data[174] = 16'b1011000000000000;
  assign in_re_table_data[175] = 16'b1011000000000000;
  assign in_re_table_data[176] = 16'b1011000000000000;
  assign in_re_table_data[177] = 16'b1011001000000000;
  assign in_re_table_data[178] = 16'b1011011000000000;
  assign in_re_table_data[179] = 16'b1011101000000000;
  assign in_re_table_data[180] = 16'b1100000000000000;
  assign in_re_table_data[181] = 16'b1100011000000000;
  assign in_re_table_data[182] = 16'b1100111000000000;
  assign in_re_table_data[183] = 16'b1101010111111111;
  assign in_re_table_data[184] = 16'b1101111000000000;
  assign in_re_table_data[185] = 16'b1110011111111111;
  assign in_re_table_data[186] = 16'b1111000111111111;
  assign in_re_table_data[187] = 16'b1111101000000000;
  assign in_re_table_data[188] = 16'b0000010111111111;
  assign in_re_table_data[189] = 16'b0000110111111111;
  assign in_re_table_data[190] = 16'b0001011111111111;
  assign in_re_table_data[191] = 16'b0010000111111111;
  assign in_re_table_data[192] = 16'b0010101000000000;
  assign in_re_table_data[193] = 16'b0011000111111111;
  assign in_re_table_data[194] = 16'b0011101000000000;
  assign in_re_table_data[195] = 16'b0100000000000000;
  assign in_re_table_data[196] = 16'b0100011000000000;
  assign in_re_table_data[197] = 16'b0100100111111111;
  assign in_re_table_data[198] = 16'b0100111000000000;
  assign in_re_table_data[199] = 16'b0101000000000000;
  assign in_re_table_data[200] = 16'b0100111111111111;
  assign in_re_table_data[201] = 16'b0101000000000000;
  assign in_re_table_data[202] = 16'b0100110111111111;
  assign in_re_table_data[203] = 16'b0100100111111111;
  assign in_re_table_data[204] = 16'b0100010111111111;
  assign in_re_table_data[205] = 16'b0100000000000000;
  assign in_re_table_data[206] = 16'b0011100111111111;
  assign in_re_table_data[207] = 16'b0011000111111111;
  assign in_re_table_data[208] = 16'b0010100111111111;
  assign in_re_table_data[209] = 16'b0010001000000000;
  assign in_re_table_data[210] = 16'b0001011111111111;
  assign in_re_table_data[211] = 16'b0000111000000000;
  assign in_re_table_data[212] = 16'b0000011000000000;
  assign in_re_table_data[213] = 16'b1111101000000000;
  assign in_re_table_data[214] = 16'b1111001000000000;
  assign in_re_table_data[215] = 16'b1110100000000000;
  assign in_re_table_data[216] = 16'b1101111000000000;
  assign in_re_table_data[217] = 16'b1101011000000000;
  assign in_re_table_data[218] = 16'b1100111000000000;
  assign in_re_table_data[219] = 16'b1100011000000000;
  assign in_re_table_data[220] = 16'b1100000000000000;
  assign in_re_table_data[221] = 16'b1011101000000000;
  assign in_re_table_data[222] = 16'b1011011000000000;
  assign in_re_table_data[223] = 16'b1011001000000000;
  assign in_re_table_data[224] = 16'b1011000000000000;
  assign in_re_table_data[225] = 16'b1011000000000000;
  assign in_re_table_data[226] = 16'b1011000000000000;
  assign in_re_table_data[227] = 16'b1011001000000000;
  assign in_re_table_data[228] = 16'b1011011000000000;
  assign in_re_table_data[229] = 16'b1011101000000000;
  assign in_re_table_data[230] = 16'b1100000000000000;
  assign in_re_table_data[231] = 16'b1100011000000000;
  assign in_re_table_data[232] = 16'b1100111000000000;
  assign in_re_table_data[233] = 16'b1101010111111111;
  assign in_re_table_data[234] = 16'b1101111000000000;
  assign in_re_table_data[235] = 16'b1110011111111111;
  assign in_re_table_data[236] = 16'b1111000111111111;
  assign in_re_table_data[237] = 16'b1111101000000000;
  assign in_re_table_data[238] = 16'b0000010111111111;
  assign in_re_table_data[239] = 16'b0000110111111111;
  assign in_re_table_data[240] = 16'b0001011111111111;
  assign in_re_table_data[241] = 16'b0010000111111111;
  assign in_re_table_data[242] = 16'b0010101000000000;
  assign in_re_table_data[243] = 16'b0011000111111111;
  assign in_re_table_data[244] = 16'b0011101000000000;
  assign in_re_table_data[245] = 16'b0100000000000000;
  assign in_re_table_data[246] = 16'b0100011000000000;
  assign in_re_table_data[247] = 16'b0100100111111111;
  assign in_re_table_data[248] = 16'b0100111000000000;
  assign in_re_table_data[249] = 16'b0101000000000000;
  assign in_re_table_data[250] = 16'b1110011000000000;
  assign in_re_table_data[251] = 16'b1110011000000000;
  assign in_re_table_data[252] = 16'b1110011111111111;
  assign in_re_table_data[253] = 16'b1110100000000000;
  assign in_re_table_data[254] = 16'b1110101000000000;
  assign in_re_table_data[255] = 16'b1110110000000000;
  assign in_re_table_data[256] = 16'b1110111000000000;
  assign in_re_table_data[257] = 16'b1111000000000000;
  assign in_re_table_data[258] = 16'b1111001000000000;
  assign in_re_table_data[259] = 16'b1111010111111111;
  assign in_re_table_data[260] = 16'b1111011111111111;
  assign in_re_table_data[261] = 16'b1111110000000000;
  assign in_re_table_data[262] = 16'b1111110111111111;
  assign in_re_table_data[263] = 16'b0000000111111111;
  assign in_re_table_data[264] = 16'b0000001111111111;
  assign in_re_table_data[265] = 16'b0000011111111111;
  assign in_re_table_data[266] = 16'b0000101000000000;
  assign in_re_table_data[267] = 16'b0000111000000000;
  assign in_re_table_data[268] = 16'b0001000000000000;
  assign in_re_table_data[269] = 16'b0001000111111111;
  assign in_re_table_data[270] = 16'b0001010000000000;
  assign in_re_table_data[271] = 16'b0001011000000000;
  assign in_re_table_data[272] = 16'b0001100000000000;
  assign in_re_table_data[273] = 16'b0001100000000000;
  assign in_re_table_data[274] = 16'b0001100111111111;
  assign in_re_table_data[275] = 16'b0001101000000000;
  assign in_re_table_data[276] = 16'b0001100111111111;
  assign in_re_table_data[277] = 16'b0001100000000000;
  assign in_re_table_data[278] = 16'b0001100000000000;
  assign in_re_table_data[279] = 16'b0001011000000000;
  assign in_re_table_data[280] = 16'b0001010000000000;
  assign in_re_table_data[281] = 16'b0001001000000000;
  assign in_re_table_data[282] = 16'b0001000000000000;
  assign in_re_table_data[283] = 16'b0000111000000000;
  assign in_re_table_data[284] = 16'b0000100111111111;
  assign in_re_table_data[285] = 16'b0000100000000000;
  assign in_re_table_data[286] = 16'b0000001111111111;
  assign in_re_table_data[287] = 16'b0000001000000000;
  assign in_re_table_data[288] = 16'b1111111000000000;
  assign in_re_table_data[289] = 16'b1111110000000000;
  assign in_re_table_data[290] = 16'b1111011111111111;
  assign in_re_table_data[291] = 16'b1111010111111111;
  assign in_re_table_data[292] = 16'b1111000111111111;
  assign in_re_table_data[293] = 16'b1111000000000000;
  assign in_re_table_data[294] = 16'b1110111000000000;
  assign in_re_table_data[295] = 16'b1110110000000000;
  assign in_re_table_data[296] = 16'b1110101000000000;
  assign in_re_table_data[297] = 16'b1110100000000000;
  assign in_re_table_data[298] = 16'b1110100000000000;
  assign in_re_table_data[299] = 16'b1110011000000000;
  assign in_re_table_data[300] = 16'b1110011000000000;
  assign in_re_table_data[301] = 16'b1110011000000000;
  assign in_re_table_data[302] = 16'b1110011111111111;
  assign in_re_table_data[303] = 16'b1110100000000000;
  assign in_re_table_data[304] = 16'b1110101000000000;
  assign in_re_table_data[305] = 16'b1110110000000000;
  assign in_re_table_data[306] = 16'b1110111000000000;
  assign in_re_table_data[307] = 16'b1111000000000000;
  assign in_re_table_data[308] = 16'b1111001000000000;
  assign in_re_table_data[309] = 16'b1111010111111111;
  assign in_re_table_data[310] = 16'b1111011111111111;
  assign in_re_table_data[311] = 16'b1111110000000000;
  assign in_re_table_data[312] = 16'b1111110111111111;
  assign in_re_table_data[313] = 16'b0000000111111111;
  assign in_re_table_data[314] = 16'b0000001111111111;
  assign in_re_table_data[315] = 16'b0000011111111111;
  assign in_re_table_data[316] = 16'b0000101000000000;
  assign in_re_table_data[317] = 16'b0000111000000000;
  assign in_re_table_data[318] = 16'b0001000000000000;
  assign in_re_table_data[319] = 16'b0001000111111111;
  assign in_re_table_data[320] = 16'b0001010000000000;
  assign in_re_table_data[321] = 16'b0001011000000000;
  assign in_re_table_data[322] = 16'b0001100000000000;
  assign in_re_table_data[323] = 16'b0001100000000000;
  assign in_re_table_data[324] = 16'b0001100111111111;
  assign in_re_table_data[325] = 16'b0001101000000000;
  assign in_re_table_data[326] = 16'b0001100111111111;
  assign in_re_table_data[327] = 16'b0001100000000000;
  assign in_re_table_data[328] = 16'b0001100000000000;
  assign in_re_table_data[329] = 16'b0001011000000000;
  assign in_re_table_data[330] = 16'b0001010000000000;
  assign in_re_table_data[331] = 16'b0001001000000000;
  assign in_re_table_data[332] = 16'b0001000000000000;
  assign in_re_table_data[333] = 16'b0000111000000000;
  assign in_re_table_data[334] = 16'b0000100111111111;
  assign in_re_table_data[335] = 16'b0000100000000000;
  assign in_re_table_data[336] = 16'b0000001111111111;
  assign in_re_table_data[337] = 16'b0000001000000000;
  assign in_re_table_data[338] = 16'b1111111000000000;
  assign in_re_table_data[339] = 16'b1111110000000000;
  assign in_re_table_data[340] = 16'b1111011111111111;
  assign in_re_table_data[341] = 16'b1111010111111111;
  assign in_re_table_data[342] = 16'b1111000111111111;
  assign in_re_table_data[343] = 16'b1111000000000000;
  assign in_re_table_data[344] = 16'b1110111000000000;
  assign in_re_table_data[345] = 16'b1110110000000000;
  assign in_re_table_data[346] = 16'b1110101000000000;
  assign in_re_table_data[347] = 16'b1110100000000000;
  assign in_re_table_data[348] = 16'b1110100000000000;
  assign in_re_table_data[349] = 16'b1110011000000000;
  assign in_re_table_data[350] = 16'b1110011000000000;
  assign in_re_table_data[351] = 16'b1110011000000000;
  assign in_re_table_data[352] = 16'b1110011111111111;
  assign in_re_table_data[353] = 16'b1110100000000000;
  assign in_re_table_data[354] = 16'b1110101000000000;
  assign in_re_table_data[355] = 16'b1110110000000000;
  assign in_re_table_data[356] = 16'b1110111000000000;
  assign in_re_table_data[357] = 16'b1111000000000000;
  assign in_re_table_data[358] = 16'b1111001000000000;
  assign in_re_table_data[359] = 16'b1111010111111111;
  assign in_re_table_data[360] = 16'b1111011111111111;
  assign in_re_table_data[361] = 16'b1111110000000000;
  assign in_re_table_data[362] = 16'b1111110111111111;
  assign in_re_table_data[363] = 16'b0000000111111111;
  assign in_re_table_data[364] = 16'b0000001111111111;
  assign in_re_table_data[365] = 16'b0000011111111111;
  assign in_re_table_data[366] = 16'b0000101000000000;
  assign in_re_table_data[367] = 16'b0000111000000000;
  assign in_re_table_data[368] = 16'b0001000000000000;
  assign in_re_table_data[369] = 16'b0001000111111111;
  assign in_re_table_data[370] = 16'b0001010000000000;
  assign in_re_table_data[371] = 16'b0001011000000000;
  assign in_re_table_data[372] = 16'b0001100000000000;
  assign in_re_table_data[373] = 16'b0001100000000000;
  assign in_re_table_data[374] = 16'b0001100111111111;
  assign in_re_table_data[375] = 16'b0001101000000000;
  assign in_re_table_data[376] = 16'b0001100111111111;
  assign in_re_table_data[377] = 16'b0001100000000000;
  assign in_re_table_data[378] = 16'b0001100000000000;
  assign in_re_table_data[379] = 16'b0001011000000000;
  assign in_re_table_data[380] = 16'b0001010000000000;
  assign in_re_table_data[381] = 16'b0001001000000000;
  assign in_re_table_data[382] = 16'b0001000000000000;
  assign in_re_table_data[383] = 16'b0000111000000000;
  assign in_re_table_data[384] = 16'b0000100111111111;
  assign in_re_table_data[385] = 16'b0000100000000000;
  assign in_re_table_data[386] = 16'b0000001111111111;
  assign in_re_table_data[387] = 16'b0000001000000000;
  assign in_re_table_data[388] = 16'b1111111000000000;
  assign in_re_table_data[389] = 16'b1111110000000000;
  assign in_re_table_data[390] = 16'b1111011111111111;
  assign in_re_table_data[391] = 16'b1111010111111111;
  assign in_re_table_data[392] = 16'b1111000111111111;
  assign in_re_table_data[393] = 16'b1111000000000000;
  assign in_re_table_data[394] = 16'b1110111000000000;
  assign in_re_table_data[395] = 16'b1110110000000000;
  assign in_re_table_data[396] = 16'b1110101000000000;
  assign in_re_table_data[397] = 16'b1110100000000000;
  assign in_re_table_data[398] = 16'b1110100000000000;
  assign in_re_table_data[399] = 16'b1110011000000000;
  assign in_re_table_data[400] = 16'b1110011000000000;
  assign in_re_table_data[401] = 16'b1110011000000000;
  assign in_re_table_data[402] = 16'b1110011111111111;
  assign in_re_table_data[403] = 16'b1110100000000000;
  assign in_re_table_data[404] = 16'b1110101000000000;
  assign in_re_table_data[405] = 16'b1110110000000000;
  assign in_re_table_data[406] = 16'b1110111000000000;
  assign in_re_table_data[407] = 16'b1111000000000000;
  assign in_re_table_data[408] = 16'b1111001000000000;
  assign in_re_table_data[409] = 16'b1111010111111111;
  assign in_re_table_data[410] = 16'b1111011111111111;
  assign in_re_table_data[411] = 16'b1111110000000000;
  assign in_re_table_data[412] = 16'b1111110111111111;
  assign in_re_table_data[413] = 16'b0000000111111111;
  assign in_re_table_data[414] = 16'b0000001111111111;
  assign in_re_table_data[415] = 16'b0000011111111111;
  assign in_re_table_data[416] = 16'b0000101000000000;
  assign in_re_table_data[417] = 16'b0000111000000000;
  assign in_re_table_data[418] = 16'b0001000000000000;
  assign in_re_table_data[419] = 16'b0001000111111111;
  assign in_re_table_data[420] = 16'b0001010000000000;
  assign in_re_table_data[421] = 16'b0001011000000000;
  assign in_re_table_data[422] = 16'b0001100000000000;
  assign in_re_table_data[423] = 16'b0001100000000000;
  assign in_re_table_data[424] = 16'b0001100111111111;
  assign in_re_table_data[425] = 16'b0001101000000000;
  assign in_re_table_data[426] = 16'b0001100111111111;
  assign in_re_table_data[427] = 16'b0001100000000000;
  assign in_re_table_data[428] = 16'b0001100000000000;
  assign in_re_table_data[429] = 16'b0001011000000000;
  assign in_re_table_data[430] = 16'b0001010000000000;
  assign in_re_table_data[431] = 16'b0001001000000000;
  assign in_re_table_data[432] = 16'b0001000000000000;
  assign in_re_table_data[433] = 16'b0000111000000000;
  assign in_re_table_data[434] = 16'b0000100111111111;
  assign in_re_table_data[435] = 16'b0000100000000000;
  assign in_re_table_data[436] = 16'b0000001111111111;
  assign in_re_table_data[437] = 16'b0000001000000000;
  assign in_re_table_data[438] = 16'b1111111000000000;
  assign in_re_table_data[439] = 16'b1111110000000000;
  assign in_re_table_data[440] = 16'b1111011111111111;
  assign in_re_table_data[441] = 16'b1111010111111111;
  assign in_re_table_data[442] = 16'b1111000111111111;
  assign in_re_table_data[443] = 16'b1111000000000000;
  assign in_re_table_data[444] = 16'b1110111000000000;
  assign in_re_table_data[445] = 16'b1110110000000000;
  assign in_re_table_data[446] = 16'b1110101000000000;
  assign in_re_table_data[447] = 16'b1110100000000000;
  assign in_re_table_data[448] = 16'b1110100000000000;
  assign in_re_table_data[449] = 16'b1110011000000000;
  assign in_re_table_data[450] = 16'b1110011000000000;
  assign in_re_table_data[451] = 16'b1110011000000000;
  assign in_re_table_data[452] = 16'b1110011111111111;
  assign in_re_table_data[453] = 16'b1110100000000000;
  assign in_re_table_data[454] = 16'b1110101000000000;
  assign in_re_table_data[455] = 16'b1110110000000000;
  assign in_re_table_data[456] = 16'b1110111000000000;
  assign in_re_table_data[457] = 16'b1111000000000000;
  assign in_re_table_data[458] = 16'b1111001000000000;
  assign in_re_table_data[459] = 16'b1111010111111111;
  assign in_re_table_data[460] = 16'b1111011111111111;
  assign in_re_table_data[461] = 16'b1111110000000000;
  assign in_re_table_data[462] = 16'b1111110111111111;
  assign in_re_table_data[463] = 16'b0000000111111111;
  assign in_re_table_data[464] = 16'b0000001111111111;
  assign in_re_table_data[465] = 16'b0000011111111111;
  assign in_re_table_data[466] = 16'b0000101000000000;
  assign in_re_table_data[467] = 16'b0000111000000000;
  assign in_re_table_data[468] = 16'b0001000000000000;
  assign in_re_table_data[469] = 16'b0001000111111111;
  assign in_re_table_data[470] = 16'b0001010000000000;
  assign in_re_table_data[471] = 16'b0001011000000000;
  assign in_re_table_data[472] = 16'b0001100000000000;
  assign in_re_table_data[473] = 16'b0001100000000000;
  assign in_re_table_data[474] = 16'b0001100111111111;
  assign in_re_table_data[475] = 16'b0001101000000000;
  assign in_re_table_data[476] = 16'b0001100111111111;
  assign in_re_table_data[477] = 16'b0001100000000000;
  assign in_re_table_data[478] = 16'b0001100000000000;
  assign in_re_table_data[479] = 16'b0001011000000000;
  assign in_re_table_data[480] = 16'b0001010000000000;
  assign in_re_table_data[481] = 16'b0001001000000000;
  assign in_re_table_data[482] = 16'b0001000000000000;
  assign in_re_table_data[483] = 16'b0000111000000000;
  assign in_re_table_data[484] = 16'b0000100111111111;
  assign in_re_table_data[485] = 16'b0000100000000000;
  assign in_re_table_data[486] = 16'b0000001111111111;
  assign in_re_table_data[487] = 16'b0000001000000000;
  assign in_re_table_data[488] = 16'b1111111000000000;
  assign in_re_table_data[489] = 16'b1111110000000000;
  assign in_re_table_data[490] = 16'b1111011111111111;
  assign in_re_table_data[491] = 16'b1111010111111111;
  assign in_re_table_data[492] = 16'b1111000111111111;
  assign in_re_table_data[493] = 16'b1111000000000000;
  assign in_re_table_data[494] = 16'b1110111000000000;
  assign in_re_table_data[495] = 16'b1110110000000000;
  assign in_re_table_data[496] = 16'b1110101000000000;
  assign in_re_table_data[497] = 16'b1110100000000000;
  assign in_re_table_data[498] = 16'b1110100000000000;
  assign in_re_table_data[499] = 16'b1110011000000000;
  assign in_re_table_data[500] = 16'b0001000111111111;
  assign in_re_table_data[501] = 16'b0001010111111111;
  assign in_re_table_data[502] = 16'b0001100111111111;
  assign in_re_table_data[503] = 16'b0001110000000000;
  assign in_re_table_data[504] = 16'b0001111000000000;
  assign in_re_table_data[505] = 16'b0010000000000000;
  assign in_re_table_data[506] = 16'b0010000111111111;
  assign in_re_table_data[507] = 16'b0010010000000000;
  assign in_re_table_data[508] = 16'b0010001111111111;
  assign in_re_table_data[509] = 16'b0010010000000000;
  assign in_re_table_data[510] = 16'b0010010000000000;
  assign in_re_table_data[511] = 16'b0010001000000000;
  assign in_re_table_data[512] = 16'b0001111111111111;
  assign in_re_table_data[513] = 16'b0001110111111111;
  assign in_re_table_data[514] = 16'b0001110000000000;
  assign in_re_table_data[515] = 16'b0001100000000000;
  assign in_re_table_data[516] = 16'b0001010000000000;
  assign in_re_table_data[517] = 16'b0000111111111111;
  assign in_re_table_data[518] = 16'b0000101111111111;
  assign in_re_table_data[519] = 16'b0000011111111111;
  assign in_re_table_data[520] = 16'b0000010000000000;
  assign in_re_table_data[521] = 16'b1111111111111111;
  assign in_re_table_data[522] = 16'b1111100111111111;
  assign in_re_table_data[523] = 16'b1111010111111111;
  assign in_re_table_data[524] = 16'b1111000111111111;
  assign in_re_table_data[525] = 16'b1110111000000000;
  assign in_re_table_data[526] = 16'b1110101000000000;
  assign in_re_table_data[527] = 16'b1110010111111111;
  assign in_re_table_data[528] = 16'b1110010000000000;
  assign in_re_table_data[529] = 16'b1110001000000000;
  assign in_re_table_data[530] = 16'b1110000000000000;
  assign in_re_table_data[531] = 16'b1101111000000000;
  assign in_re_table_data[532] = 16'b1101110000000000;
  assign in_re_table_data[533] = 16'b1101110000000000;
  assign in_re_table_data[534] = 16'b1101101111111111;
  assign in_re_table_data[535] = 16'b1101101111111111;
  assign in_re_table_data[536] = 16'b1101111000000000;
  assign in_re_table_data[537] = 16'b1110000000000000;
  assign in_re_table_data[538] = 16'b1110001000000000;
  assign in_re_table_data[539] = 16'b1110010000000000;
  assign in_re_table_data[540] = 16'b1110100000000000;
  assign in_re_table_data[541] = 16'b1110110000000000;
  assign in_re_table_data[542] = 16'b1111000000000000;
  assign in_re_table_data[543] = 16'b1111010000000000;
  assign in_re_table_data[544] = 16'b1111100000000000;
  assign in_re_table_data[545] = 16'b1111101111111111;
  assign in_re_table_data[546] = 16'b0000000000000000;
  assign in_re_table_data[547] = 16'b0000011000000000;
  assign in_re_table_data[548] = 16'b0000101000000000;
  assign in_re_table_data[549] = 16'b0000111000000000;
  assign in_re_table_data[550] = 16'b0001000111111111;
  assign in_re_table_data[551] = 16'b0001010111111111;
  assign in_re_table_data[552] = 16'b0001100111111111;
  assign in_re_table_data[553] = 16'b0001110000000000;
  assign in_re_table_data[554] = 16'b0001111000000000;
  assign in_re_table_data[555] = 16'b0010000000000000;
  assign in_re_table_data[556] = 16'b0010000111111111;
  assign in_re_table_data[557] = 16'b0010010000000000;
  assign in_re_table_data[558] = 16'b0010001111111111;
  assign in_re_table_data[559] = 16'b0010010000000000;
  assign in_re_table_data[560] = 16'b0010010000000000;
  assign in_re_table_data[561] = 16'b0010001000000000;
  assign in_re_table_data[562] = 16'b0001111111111111;
  assign in_re_table_data[563] = 16'b0001110111111111;
  assign in_re_table_data[564] = 16'b0001110000000000;
  assign in_re_table_data[565] = 16'b0001100000000000;
  assign in_re_table_data[566] = 16'b0001010000000000;
  assign in_re_table_data[567] = 16'b0000111111111111;
  assign in_re_table_data[568] = 16'b0000101111111111;
  assign in_re_table_data[569] = 16'b0000011111111111;
  assign in_re_table_data[570] = 16'b0000010000000000;
  assign in_re_table_data[571] = 16'b1111111111111111;
  assign in_re_table_data[572] = 16'b1111100111111111;
  assign in_re_table_data[573] = 16'b1111010111111111;
  assign in_re_table_data[574] = 16'b1111000111111111;
  assign in_re_table_data[575] = 16'b1110111000000000;
  assign in_re_table_data[576] = 16'b1110101000000000;
  assign in_re_table_data[577] = 16'b1110010111111111;
  assign in_re_table_data[578] = 16'b1110010000000000;
  assign in_re_table_data[579] = 16'b1110001000000000;
  assign in_re_table_data[580] = 16'b1110000000000000;
  assign in_re_table_data[581] = 16'b1101111000000000;
  assign in_re_table_data[582] = 16'b1101110000000000;
  assign in_re_table_data[583] = 16'b1101110000000000;
  assign in_re_table_data[584] = 16'b1101101111111111;
  assign in_re_table_data[585] = 16'b1101101111111111;
  assign in_re_table_data[586] = 16'b1101111000000000;
  assign in_re_table_data[587] = 16'b1110000000000000;
  assign in_re_table_data[588] = 16'b1110001000000000;
  assign in_re_table_data[589] = 16'b1110010000000000;
  assign in_re_table_data[590] = 16'b1110100000000000;
  assign in_re_table_data[591] = 16'b1110110000000000;
  assign in_re_table_data[592] = 16'b1111000000000000;
  assign in_re_table_data[593] = 16'b1111010000000000;
  assign in_re_table_data[594] = 16'b1111100000000000;
  assign in_re_table_data[595] = 16'b1111101111111111;
  assign in_re_table_data[596] = 16'b0000000000000000;
  assign in_re_table_data[597] = 16'b0000011000000000;
  assign in_re_table_data[598] = 16'b0000101000000000;
  assign in_re_table_data[599] = 16'b0000111000000000;
  assign in_re_table_data[600] = 16'b0001000111111111;
  assign in_re_table_data[601] = 16'b0001010111111111;
  assign in_re_table_data[602] = 16'b0001100111111111;
  assign in_re_table_data[603] = 16'b0001110000000000;
  assign in_re_table_data[604] = 16'b0001111000000000;
  assign in_re_table_data[605] = 16'b0010000000000000;
  assign in_re_table_data[606] = 16'b0010000111111111;
  assign in_re_table_data[607] = 16'b0010010000000000;
  assign in_re_table_data[608] = 16'b0010001111111111;
  assign in_re_table_data[609] = 16'b0010010000000000;
  assign in_re_table_data[610] = 16'b0010010000000000;
  assign in_re_table_data[611] = 16'b0010001000000000;
  assign in_re_table_data[612] = 16'b0001111111111111;
  assign in_re_table_data[613] = 16'b0001110111111111;
  assign in_re_table_data[614] = 16'b0001110000000000;
  assign in_re_table_data[615] = 16'b0001100000000000;
  assign in_re_table_data[616] = 16'b0001010000000000;
  assign in_re_table_data[617] = 16'b0000111111111111;
  assign in_re_table_data[618] = 16'b0000101111111111;
  assign in_re_table_data[619] = 16'b0000011111111111;
  assign in_re_table_data[620] = 16'b0000010000000000;
  assign in_re_table_data[621] = 16'b1111111111111111;
  assign in_re_table_data[622] = 16'b1111100111111111;
  assign in_re_table_data[623] = 16'b1111010111111111;
  assign in_re_table_data[624] = 16'b1111000111111111;
  assign in_re_table_data[625] = 16'b1110111000000000;
  assign in_re_table_data[626] = 16'b1110101000000000;
  assign in_re_table_data[627] = 16'b1110010111111111;
  assign in_re_table_data[628] = 16'b1110010000000000;
  assign in_re_table_data[629] = 16'b1110001000000000;
  assign in_re_table_data[630] = 16'b1110000000000000;
  assign in_re_table_data[631] = 16'b1101111000000000;
  assign in_re_table_data[632] = 16'b1101110000000000;
  assign in_re_table_data[633] = 16'b1101110000000000;
  assign in_re_table_data[634] = 16'b1101101111111111;
  assign in_re_table_data[635] = 16'b1101101111111111;
  assign in_re_table_data[636] = 16'b1101111000000000;
  assign in_re_table_data[637] = 16'b1110000000000000;
  assign in_re_table_data[638] = 16'b1110001000000000;
  assign in_re_table_data[639] = 16'b1110010000000000;
  assign in_re_table_data[640] = 16'b1110100000000000;
  assign in_re_table_data[641] = 16'b1110110000000000;
  assign in_re_table_data[642] = 16'b1111000000000000;
  assign in_re_table_data[643] = 16'b1111010000000000;
  assign in_re_table_data[644] = 16'b1111100000000000;
  assign in_re_table_data[645] = 16'b1111101111111111;
  assign in_re_table_data[646] = 16'b0000000000000000;
  assign in_re_table_data[647] = 16'b0000011000000000;
  assign in_re_table_data[648] = 16'b0000101000000000;
  assign in_re_table_data[649] = 16'b0000111000000000;
  assign in_re_table_data[650] = 16'b0001000111111111;
  assign in_re_table_data[651] = 16'b0001010111111111;
  assign in_re_table_data[652] = 16'b0001100111111111;
  assign in_re_table_data[653] = 16'b0001110000000000;
  assign in_re_table_data[654] = 16'b0001111000000000;
  assign in_re_table_data[655] = 16'b0010000000000000;
  assign in_re_table_data[656] = 16'b0010000111111111;
  assign in_re_table_data[657] = 16'b0010010000000000;
  assign in_re_table_data[658] = 16'b0010001111111111;
  assign in_re_table_data[659] = 16'b0010010000000000;
  assign in_re_table_data[660] = 16'b0010010000000000;
  assign in_re_table_data[661] = 16'b0010001000000000;
  assign in_re_table_data[662] = 16'b0001111111111111;
  assign in_re_table_data[663] = 16'b0001110111111111;
  assign in_re_table_data[664] = 16'b0001110000000000;
  assign in_re_table_data[665] = 16'b0001100000000000;
  assign in_re_table_data[666] = 16'b0001010000000000;
  assign in_re_table_data[667] = 16'b0000111111111111;
  assign in_re_table_data[668] = 16'b0000101111111111;
  assign in_re_table_data[669] = 16'b0000011111111111;
  assign in_re_table_data[670] = 16'b0000010000000000;
  assign in_re_table_data[671] = 16'b1111111111111111;
  assign in_re_table_data[672] = 16'b1111100111111111;
  assign in_re_table_data[673] = 16'b1111010111111111;
  assign in_re_table_data[674] = 16'b1111000111111111;
  assign in_re_table_data[675] = 16'b1110111000000000;
  assign in_re_table_data[676] = 16'b1110101000000000;
  assign in_re_table_data[677] = 16'b1110010111111111;
  assign in_re_table_data[678] = 16'b1110010000000000;
  assign in_re_table_data[679] = 16'b1110001000000000;
  assign in_re_table_data[680] = 16'b1110000000000000;
  assign in_re_table_data[681] = 16'b1101111000000000;
  assign in_re_table_data[682] = 16'b1101110000000000;
  assign in_re_table_data[683] = 16'b1101110000000000;
  assign in_re_table_data[684] = 16'b1101101111111111;
  assign in_re_table_data[685] = 16'b1101101111111111;
  assign in_re_table_data[686] = 16'b1101111000000000;
  assign in_re_table_data[687] = 16'b1110000000000000;
  assign in_re_table_data[688] = 16'b1110001000000000;
  assign in_re_table_data[689] = 16'b1110010000000000;
  assign in_re_table_data[690] = 16'b1110100000000000;
  assign in_re_table_data[691] = 16'b1110110000000000;
  assign in_re_table_data[692] = 16'b1111000000000000;
  assign in_re_table_data[693] = 16'b1111010000000000;
  assign in_re_table_data[694] = 16'b1111100000000000;
  assign in_re_table_data[695] = 16'b1111101111111111;
  assign in_re_table_data[696] = 16'b0000000000000000;
  assign in_re_table_data[697] = 16'b0000011000000000;
  assign in_re_table_data[698] = 16'b0000101000000000;
  assign in_re_table_data[699] = 16'b0000111000000000;
  assign in_re_table_data[700] = 16'b0001000111111111;
  assign in_re_table_data[701] = 16'b0001010111111111;
  assign in_re_table_data[702] = 16'b0001100111111111;
  assign in_re_table_data[703] = 16'b0001110000000000;
  assign in_re_table_data[704] = 16'b0001111000000000;
  assign in_re_table_data[705] = 16'b0010000000000000;
  assign in_re_table_data[706] = 16'b0010000111111111;
  assign in_re_table_data[707] = 16'b0010010000000000;
  assign in_re_table_data[708] = 16'b0010001111111111;
  assign in_re_table_data[709] = 16'b0010010000000000;
  assign in_re_table_data[710] = 16'b0010010000000000;
  assign in_re_table_data[711] = 16'b0010001000000000;
  assign in_re_table_data[712] = 16'b0001111111111111;
  assign in_re_table_data[713] = 16'b0001110111111111;
  assign in_re_table_data[714] = 16'b0001110000000000;
  assign in_re_table_data[715] = 16'b0001100000000000;
  assign in_re_table_data[716] = 16'b0001010000000000;
  assign in_re_table_data[717] = 16'b0000111111111111;
  assign in_re_table_data[718] = 16'b0000101111111111;
  assign in_re_table_data[719] = 16'b0000011111111111;
  assign in_re_table_data[720] = 16'b0000010000000000;
  assign in_re_table_data[721] = 16'b1111111111111111;
  assign in_re_table_data[722] = 16'b1111100111111111;
  assign in_re_table_data[723] = 16'b1111010111111111;
  assign in_re_table_data[724] = 16'b1111000111111111;
  assign in_re_table_data[725] = 16'b1110111000000000;
  assign in_re_table_data[726] = 16'b1110101000000000;
  assign in_re_table_data[727] = 16'b1110010111111111;
  assign in_re_table_data[728] = 16'b1110010000000000;
  assign in_re_table_data[729] = 16'b1110001000000000;
  assign in_re_table_data[730] = 16'b1110000000000000;
  assign in_re_table_data[731] = 16'b1101111000000000;
  assign in_re_table_data[732] = 16'b1101110000000000;
  assign in_re_table_data[733] = 16'b1101110000000000;
  assign in_re_table_data[734] = 16'b1101101111111111;
  assign in_re_table_data[735] = 16'b1101101111111111;
  assign in_re_table_data[736] = 16'b1101111000000000;
  assign in_re_table_data[737] = 16'b1110000000000000;
  assign in_re_table_data[738] = 16'b1110001000000000;
  assign in_re_table_data[739] = 16'b1110010000000000;
  assign in_re_table_data[740] = 16'b1110100000000000;
  assign in_re_table_data[741] = 16'b1110110000000000;
  assign in_re_table_data[742] = 16'b1111000000000000;
  assign in_re_table_data[743] = 16'b1111010000000000;
  assign in_re_table_data[744] = 16'b1111100000000000;
  assign in_re_table_data[745] = 16'b1111101111111111;
  assign in_re_table_data[746] = 16'b0000000000000000;
  assign in_re_table_data[747] = 16'b0000011000000000;
  assign in_re_table_data[748] = 16'b0000101000000000;
  assign in_re_table_data[749] = 16'b0000111000000000;
  assign in_re_table_data[750] = 16'b0000001000000000;
  assign in_re_table_data[751] = 16'b0000000111111111;
  assign in_re_table_data[752] = 16'b0000000111111111;
  assign in_re_table_data[753] = 16'b0000001000000000;
  assign in_re_table_data[754] = 16'b0000000111111111;
  assign in_re_table_data[755] = 16'b0000001000000000;
  assign in_re_table_data[756] = 16'b0000001000000000;
  assign in_re_table_data[757] = 16'b1111111111111111;
  assign in_re_table_data[758] = 16'b0000000000000000;
  assign in_re_table_data[759] = 16'b1111111111111111;
  assign in_re_table_data[760] = 16'b1111111111111111;
  assign in_re_table_data[761] = 16'b0000000000000000;
  assign in_re_table_data[762] = 16'b1111111000000000;
  assign in_re_table_data[763] = 16'b1111111000000000;
  assign in_re_table_data[764] = 16'b1111111000000000;
  assign in_re_table_data[765] = 16'b1111111000000000;
  assign in_re_table_data[766] = 16'b1111111000000000;
  assign in_re_table_data[767] = 16'b1111111000000000;
  assign in_re_table_data[768] = 16'b1111111000000000;
  assign in_re_table_data[769] = 16'b1111111000000000;
  assign in_re_table_data[770] = 16'b1111110000000000;
  assign in_re_table_data[771] = 16'b1111110000000000;
  assign in_re_table_data[772] = 16'b1111110000000000;
  assign in_re_table_data[773] = 16'b1111110000000000;
  assign in_re_table_data[774] = 16'b1111110000000000;
  assign in_re_table_data[775] = 16'b1111110111111111;
  assign in_re_table_data[776] = 16'b1111111000000000;
  assign in_re_table_data[777] = 16'b1111111000000000;
  assign in_re_table_data[778] = 16'b1111110111111111;
  assign in_re_table_data[779] = 16'b1111111000000000;
  assign in_re_table_data[780] = 16'b1111111000000000;
  assign in_re_table_data[781] = 16'b1111110111111111;
  assign in_re_table_data[782] = 16'b1111111111111111;
  assign in_re_table_data[783] = 16'b1111111111111111;
  assign in_re_table_data[784] = 16'b0000000000000000;
  assign in_re_table_data[785] = 16'b1111111111111111;
  assign in_re_table_data[786] = 16'b1111111111111111;
  assign in_re_table_data[787] = 16'b0000001000000000;
  assign in_re_table_data[788] = 16'b0000000111111111;
  assign in_re_table_data[789] = 16'b0000001000000000;
  assign in_re_table_data[790] = 16'b0000001000000000;
  assign in_re_table_data[791] = 16'b0000000111111111;
  assign in_re_table_data[792] = 16'b0000001000000000;
  assign in_re_table_data[793] = 16'b0000001000000000;
  assign in_re_table_data[794] = 16'b0000000111111111;
  assign in_re_table_data[795] = 16'b0000010000000000;
  assign in_re_table_data[796] = 16'b0000001111111111;
  assign in_re_table_data[797] = 16'b0000001111111111;
  assign in_re_table_data[798] = 16'b0000010000000000;
  assign in_re_table_data[799] = 16'b0000001111111111;
  assign in_re_table_data[800] = 16'b0000001000000000;
  assign in_re_table_data[801] = 16'b0000000111111111;
  assign in_re_table_data[802] = 16'b0000000111111111;
  assign in_re_table_data[803] = 16'b0000001000000000;
  assign in_re_table_data[804] = 16'b0000000111111111;
  assign in_re_table_data[805] = 16'b0000001000000000;
  assign in_re_table_data[806] = 16'b0000001000000000;
  assign in_re_table_data[807] = 16'b1111111111111111;
  assign in_re_table_data[808] = 16'b0000000000000000;
  assign in_re_table_data[809] = 16'b1111111111111111;
  assign in_re_table_data[810] = 16'b1111111111111111;
  assign in_re_table_data[811] = 16'b0000000000000000;
  assign in_re_table_data[812] = 16'b1111111000000000;
  assign in_re_table_data[813] = 16'b1111111000000000;
  assign in_re_table_data[814] = 16'b1111111000000000;
  assign in_re_table_data[815] = 16'b1111111000000000;
  assign in_re_table_data[816] = 16'b1111111000000000;
  assign in_re_table_data[817] = 16'b1111111000000000;
  assign in_re_table_data[818] = 16'b1111111000000000;
  assign in_re_table_data[819] = 16'b1111111000000000;
  assign in_re_table_data[820] = 16'b1111110000000000;
  assign in_re_table_data[821] = 16'b1111110000000000;
  assign in_re_table_data[822] = 16'b1111110000000000;
  assign in_re_table_data[823] = 16'b1111110000000000;
  assign in_re_table_data[824] = 16'b1111110000000000;
  assign in_re_table_data[825] = 16'b1111110111111111;
  assign in_re_table_data[826] = 16'b1111111000000000;
  assign in_re_table_data[827] = 16'b1111111000000000;
  assign in_re_table_data[828] = 16'b1111110111111111;
  assign in_re_table_data[829] = 16'b1111111000000000;
  assign in_re_table_data[830] = 16'b1111111000000000;
  assign in_re_table_data[831] = 16'b1111110111111111;
  assign in_re_table_data[832] = 16'b1111111111111111;
  assign in_re_table_data[833] = 16'b1111111111111111;
  assign in_re_table_data[834] = 16'b0000000000000000;
  assign in_re_table_data[835] = 16'b1111111111111111;
  assign in_re_table_data[836] = 16'b1111111111111111;
  assign in_re_table_data[837] = 16'b0000001000000000;
  assign in_re_table_data[838] = 16'b0000000111111111;
  assign in_re_table_data[839] = 16'b0000001000000000;
  assign in_re_table_data[840] = 16'b0000001000000000;
  assign in_re_table_data[841] = 16'b0000000111111111;
  assign in_re_table_data[842] = 16'b0000001000000000;
  assign in_re_table_data[843] = 16'b0000001000000000;
  assign in_re_table_data[844] = 16'b0000000111111111;
  assign in_re_table_data[845] = 16'b0000010000000000;
  assign in_re_table_data[846] = 16'b0000001111111111;
  assign in_re_table_data[847] = 16'b0000001111111111;
  assign in_re_table_data[848] = 16'b0000010000000000;
  assign in_re_table_data[849] = 16'b0000001111111111;
  assign in_re_table_data[850] = 16'b0000001000000000;
  assign in_re_table_data[851] = 16'b0000000111111111;
  assign in_re_table_data[852] = 16'b0000000111111111;
  assign in_re_table_data[853] = 16'b0000001000000000;
  assign in_re_table_data[854] = 16'b0000000111111111;
  assign in_re_table_data[855] = 16'b0000001000000000;
  assign in_re_table_data[856] = 16'b0000001000000000;
  assign in_re_table_data[857] = 16'b1111111111111111;
  assign in_re_table_data[858] = 16'b0000000000000000;
  assign in_re_table_data[859] = 16'b1111111111111111;
  assign in_re_table_data[860] = 16'b1111111111111111;
  assign in_re_table_data[861] = 16'b0000000000000000;
  assign in_re_table_data[862] = 16'b1111111000000000;
  assign in_re_table_data[863] = 16'b1111111000000000;
  assign in_re_table_data[864] = 16'b1111111000000000;
  assign in_re_table_data[865] = 16'b1111111000000000;
  assign in_re_table_data[866] = 16'b1111111000000000;
  assign in_re_table_data[867] = 16'b1111111000000000;
  assign in_re_table_data[868] = 16'b1111111000000000;
  assign in_re_table_data[869] = 16'b1111111000000000;
  assign in_re_table_data[870] = 16'b1111110000000000;
  assign in_re_table_data[871] = 16'b1111110000000000;
  assign in_re_table_data[872] = 16'b1111110000000000;
  assign in_re_table_data[873] = 16'b1111110000000000;
  assign in_re_table_data[874] = 16'b1111110000000000;
  assign in_re_table_data[875] = 16'b1111110111111111;
  assign in_re_table_data[876] = 16'b1111111000000000;
  assign in_re_table_data[877] = 16'b1111111000000000;
  assign in_re_table_data[878] = 16'b1111110111111111;
  assign in_re_table_data[879] = 16'b1111111000000000;
  assign in_re_table_data[880] = 16'b1111111000000000;
  assign in_re_table_data[881] = 16'b1111110111111111;
  assign in_re_table_data[882] = 16'b1111111111111111;
  assign in_re_table_data[883] = 16'b1111111111111111;
  assign in_re_table_data[884] = 16'b0000000000000000;
  assign in_re_table_data[885] = 16'b1111111111111111;
  assign in_re_table_data[886] = 16'b1111111111111111;
  assign in_re_table_data[887] = 16'b0000001000000000;
  assign in_re_table_data[888] = 16'b0000000111111111;
  assign in_re_table_data[889] = 16'b0000001000000000;
  assign in_re_table_data[890] = 16'b0000001000000000;
  assign in_re_table_data[891] = 16'b0000000111111111;
  assign in_re_table_data[892] = 16'b0000001000000000;
  assign in_re_table_data[893] = 16'b0000001000000000;
  assign in_re_table_data[894] = 16'b0000000111111111;
  assign in_re_table_data[895] = 16'b0000010000000000;
  assign in_re_table_data[896] = 16'b0000001111111111;
  assign in_re_table_data[897] = 16'b0000001111111111;
  assign in_re_table_data[898] = 16'b0000010000000000;
  assign in_re_table_data[899] = 16'b0000001111111111;
  assign in_re_table_data[900] = 16'b0000001000000000;
  assign in_re_table_data[901] = 16'b0000000111111111;
  assign in_re_table_data[902] = 16'b0000000111111111;
  assign in_re_table_data[903] = 16'b0000001000000000;
  assign in_re_table_data[904] = 16'b0000000111111111;
  assign in_re_table_data[905] = 16'b0000001000000000;
  assign in_re_table_data[906] = 16'b0000001000000000;
  assign in_re_table_data[907] = 16'b1111111111111111;
  assign in_re_table_data[908] = 16'b0000000000000000;
  assign in_re_table_data[909] = 16'b1111111111111111;
  assign in_re_table_data[910] = 16'b1111111111111111;
  assign in_re_table_data[911] = 16'b0000000000000000;
  assign in_re_table_data[912] = 16'b1111111000000000;
  assign in_re_table_data[913] = 16'b1111111000000000;
  assign in_re_table_data[914] = 16'b1111111000000000;
  assign in_re_table_data[915] = 16'b1111111000000000;
  assign in_re_table_data[916] = 16'b1111111000000000;
  assign in_re_table_data[917] = 16'b1111111000000000;
  assign in_re_table_data[918] = 16'b1111111000000000;
  assign in_re_table_data[919] = 16'b1111111000000000;
  assign in_re_table_data[920] = 16'b1111110000000000;
  assign in_re_table_data[921] = 16'b1111110000000000;
  assign in_re_table_data[922] = 16'b1111110000000000;
  assign in_re_table_data[923] = 16'b1111110000000000;
  assign in_re_table_data[924] = 16'b1111110000000000;
  assign in_re_table_data[925] = 16'b1111110111111111;
  assign in_re_table_data[926] = 16'b1111111000000000;
  assign in_re_table_data[927] = 16'b1111111000000000;
  assign in_re_table_data[928] = 16'b1111110111111111;
  assign in_re_table_data[929] = 16'b1111111000000000;
  assign in_re_table_data[930] = 16'b1111111000000000;
  assign in_re_table_data[931] = 16'b1111110111111111;
  assign in_re_table_data[932] = 16'b1111111111111111;
  assign in_re_table_data[933] = 16'b1111111111111111;
  assign in_re_table_data[934] = 16'b0000000000000000;
  assign in_re_table_data[935] = 16'b1111111111111111;
  assign in_re_table_data[936] = 16'b1111111111111111;
  assign in_re_table_data[937] = 16'b0000001000000000;
  assign in_re_table_data[938] = 16'b0000000111111111;
  assign in_re_table_data[939] = 16'b0000001000000000;
  assign in_re_table_data[940] = 16'b0000001000000000;
  assign in_re_table_data[941] = 16'b0000000111111111;
  assign in_re_table_data[942] = 16'b0000001000000000;
  assign in_re_table_data[943] = 16'b0000001000000000;
  assign in_re_table_data[944] = 16'b0000000111111111;
  assign in_re_table_data[945] = 16'b0000010000000000;
  assign in_re_table_data[946] = 16'b0000001111111111;
  assign in_re_table_data[947] = 16'b0000001111111111;
  assign in_re_table_data[948] = 16'b0000010000000000;
  assign in_re_table_data[949] = 16'b0000001111111111;
  assign in_re_table_data[950] = 16'b0000001000000000;
  assign in_re_table_data[951] = 16'b0000000111111111;
  assign in_re_table_data[952] = 16'b0000000111111111;
  assign in_re_table_data[953] = 16'b0000001000000000;
  assign in_re_table_data[954] = 16'b0000000111111111;
  assign in_re_table_data[955] = 16'b0000001000000000;
  assign in_re_table_data[956] = 16'b0000001000000000;
  assign in_re_table_data[957] = 16'b1111111111111111;
  assign in_re_table_data[958] = 16'b0000000000000000;
  assign in_re_table_data[959] = 16'b1111111111111111;
  assign in_re_table_data[960] = 16'b1111111111111111;
  assign in_re_table_data[961] = 16'b0000000000000000;
  assign in_re_table_data[962] = 16'b1111111000000000;
  assign in_re_table_data[963] = 16'b1111111000000000;
  assign in_re_table_data[964] = 16'b1111111000000000;
  assign in_re_table_data[965] = 16'b1111111000000000;
  assign in_re_table_data[966] = 16'b1111111000000000;
  assign in_re_table_data[967] = 16'b1111111000000000;
  assign in_re_table_data[968] = 16'b1111111000000000;
  assign in_re_table_data[969] = 16'b1111111000000000;
  assign in_re_table_data[970] = 16'b1111110000000000;
  assign in_re_table_data[971] = 16'b1111110000000000;
  assign in_re_table_data[972] = 16'b1111110000000000;
  assign in_re_table_data[973] = 16'b1111110000000000;
  assign in_re_table_data[974] = 16'b1111110000000000;
  assign in_re_table_data[975] = 16'b1111110111111111;
  assign in_re_table_data[976] = 16'b1111111000000000;
  assign in_re_table_data[977] = 16'b1111111000000000;
  assign in_re_table_data[978] = 16'b1111110111111111;
  assign in_re_table_data[979] = 16'b1111111000000000;
  assign in_re_table_data[980] = 16'b1111111000000000;
  assign in_re_table_data[981] = 16'b1111110111111111;
  assign in_re_table_data[982] = 16'b1111111111111111;
  assign in_re_table_data[983] = 16'b1111111111111111;
  assign in_re_table_data[984] = 16'b0000000000000000;
  assign in_re_table_data[985] = 16'b1111111111111111;
  assign in_re_table_data[986] = 16'b1111111111111111;
  assign in_re_table_data[987] = 16'b0000001000000000;
  assign in_re_table_data[988] = 16'b0000000111111111;
  assign in_re_table_data[989] = 16'b0000001000000000;
  assign in_re_table_data[990] = 16'b0000001000000000;
  assign in_re_table_data[991] = 16'b0000000111111111;
  assign in_re_table_data[992] = 16'b0000001000000000;
  assign in_re_table_data[993] = 16'b0000001000000000;
  assign in_re_table_data[994] = 16'b0000000111111111;
  assign in_re_table_data[995] = 16'b0000010000000000;
  assign in_re_table_data[996] = 16'b0000001111111111;
  assign in_re_table_data[997] = 16'b0000001111111111;
  assign in_re_table_data[998] = 16'b0000010000000000;
  assign in_re_table_data[999] = 16'b0000001111111111;
  assign in_re_table_data[1000] = 16'b1111111111111111;
  assign in_re_1 = in_re_table_data[Data_Type_Conversion1_out1_addr];



  assign rawData_in_re = in_re_1;



  // holdData reg for Data_Type_Conversion1_out1
  always @(posedge clk)
    begin : stimuli_Data_Type_Conversion1_out1_2
      if (reset_x) begin
        holdData_in_re <= 16'bx;
      end
      else begin
        holdData_in_re <= rawData_in_re;
      end
    end

  always @(rawData_in_re or rdEnb)
    begin : stimuli_Data_Type_Conversion1_out1_3
      if (rdEnb == 1'b0) begin
        in_re_offset <= holdData_in_re;
      end
      else begin
        in_re_offset <= rawData_in_re;
      end
    end

  assign #2 in_re_2 = in_re_offset;

  assign snkDonen =  ~ snkDone;



  assign resetn =  ~ reset_x;



  assign tb_enb = resetn & snkDonen;



  // Delay inside enable generation: register depth 1
  always @(posedge clk)
    begin : u_enable_delay
      if (reset_x) begin
        tb_enb_delay <= 0;
      end
      else begin
        tb_enb_delay <= tb_enb;
      end
    end

  assign rdEnb = (snkDone == 1'b0 ? tb_enb_delay :
              1'b0);



  assign #2 clk_enable = rdEnb;

  initial
    begin : reset_x_gen
      reset_x <= 1'b1;
      # (20);
      @ (posedge clk)
      # (2);
      reset_x <= 1'b0;
    end

  always 
    begin : clk_gen
      clk <= 1'b1;
      # (5);
      clk <= 1'b0;
      # (5);
      if (snkDone == 1'b1) begin
        clk <= 1'b1;
        # (5);
        clk <= 1'b0;
        # (5);
        $stop;
      end
    end

  simulink_functio u_simulink_functio (.clk(clk),
                                       .reset_x(reset_x),
                                       .clk_enable(clk_enable),
                                       .in_re(in_re_2),  // sfix16_En14
                                       .in_im(in_im_2),  // sfix16_En14
                                      // .clk_enable(clk_enable),
                                       .magnitude(magnitude),  // ufix16_En14
                                       .alpha_arctangen(alpha_arctangen)  // sfix8_En5
                                       );

  assign magnitude_enb = clk_enable & magnitude_active;



  // Count limited, Unsigned Counter
  //  initial value   = 0
  //  step value      = 1
  //  count to value  = 1000
  always @(posedge clk)
    begin : c_2_process
      if (reset_x == 1'b1) begin
        magnitude_addr <= 10'b0000000000;
      end
      else begin
        if (magnitude_enb) begin
          if (magnitude_addr >= 10'b1111101000) begin
            magnitude_addr <= 10'b0000000000;
          end
          else begin
            magnitude_addr <= magnitude_addr + 10'b0000000001;
          end
        end
      end
    end



  assign magnitude_lastAddr = magnitude_addr >= 10'b1111101000;



  assign magnitude_done = magnitude_lastAddr & resetn;



  // Delay to allow last sim cycle to complete
  always @(posedge clk)
    begin : checkDone_1
      if (reset_x) begin
        check1_done <= 0;
      end
      else begin
        if (magnitude_done_enb) begin
          check1_done <= magnitude_done;
        end
      end
    end

  assign snkDone = check1_done & check2_done;



  // Data source for magnitude_expected
  assign magnitude_expected_table_data[0] = 16'b0000000000000000;
  assign magnitude_expected_table_data[1] = 16'b0000000000000000;
  assign magnitude_expected_table_data[2] = 16'b0000000000000000;
  assign magnitude_expected_table_data[3] = 16'b0000000000000000;
  assign magnitude_expected_table_data[4] = 16'b0000000000000000;
  assign magnitude_expected_table_data[5] = 16'b0000000000000000;
  assign magnitude_expected_table_data[6] = 16'b0000000000000000;
  assign magnitude_expected_table_data[7] = 16'b0000000000000000;
  assign magnitude_expected_table_data[8] = 16'b0000000000000000;
  assign magnitude_expected_table_data[9] = 16'b0000000000000000;
  assign magnitude_expected_table_data[10] = 16'b0000000000000000;
  assign magnitude_expected_table_data[11] = 16'b0000000000000000;
  assign magnitude_expected_table_data[12] = 16'b0000000000000000;
  assign magnitude_expected_table_data[13] = 16'b0000000000000000;
  assign magnitude_expected_table_data[14] = 16'b0000000000000000;
  assign magnitude_expected_table_data[15] = 16'b0000000000000000;
  assign magnitude_expected_table_data[16] = 16'b0000000000000000;
  assign magnitude_expected_table_data[17] = 16'b0000000000000000;
  assign magnitude_expected_table_data[18] = 16'b0000000000000000;
  assign magnitude_expected_table_data[19] = 16'b0000000000000000;
  assign magnitude_expected_table_data[20] = 16'b0000000000000000;
  assign magnitude_expected_table_data[21] = 16'b0000000000000000;
  assign magnitude_expected_table_data[22] = 16'b0000000000000000;
  assign magnitude_expected_table_data[23] = 16'b0000000000000000;
  assign magnitude_expected_table_data[24] = 16'b0000000000000000;
  assign magnitude_expected_table_data[25] = 16'b0000000000000000;
  assign magnitude_expected_table_data[26] = 16'b0100111101000000;
  assign magnitude_expected_table_data[27] = 16'b0101000100110000;
  assign magnitude_expected_table_data[28] = 16'b0101000101100000;
  assign magnitude_expected_table_data[29] = 16'b0100111100110000;
  assign magnitude_expected_table_data[30] = 16'b0101000011000000;
  assign magnitude_expected_table_data[31] = 16'b0101000001010000;
  assign magnitude_expected_table_data[32] = 16'b0100111110010000;
  assign magnitude_expected_table_data[33] = 16'b0101000000000000;
  assign magnitude_expected_table_data[34] = 16'b0100111111010000;
  assign magnitude_expected_table_data[35] = 16'b0100111101100000;
  assign magnitude_expected_table_data[36] = 16'b0101000001100000;
  assign magnitude_expected_table_data[37] = 16'b0100111011110000;
  assign magnitude_expected_table_data[38] = 16'b0100111111010000;
  assign magnitude_expected_table_data[39] = 16'b0100111111010000;
  assign magnitude_expected_table_data[40] = 16'b0100111011110000;
  assign magnitude_expected_table_data[41] = 16'b0101000001100000;
  assign magnitude_expected_table_data[42] = 16'b0100111101100000;
  assign magnitude_expected_table_data[43] = 16'b0100111111010000;
  assign magnitude_expected_table_data[44] = 16'b0101000000000000;
  assign magnitude_expected_table_data[45] = 16'b0100111110010000;
  assign magnitude_expected_table_data[46] = 16'b0101000001010000;
  assign magnitude_expected_table_data[47] = 16'b0101000011000000;
  assign magnitude_expected_table_data[48] = 16'b0100111100110000;
  assign magnitude_expected_table_data[49] = 16'b0101000101100000;
  assign magnitude_expected_table_data[50] = 16'b0101000100110000;
  assign magnitude_expected_table_data[51] = 16'b0100111101000000;
  assign magnitude_expected_table_data[52] = 16'b0101000100110000;
  assign magnitude_expected_table_data[53] = 16'b0101000101100000;
  assign magnitude_expected_table_data[54] = 16'b0100111100110000;
  assign magnitude_expected_table_data[55] = 16'b0101000011000000;
  assign magnitude_expected_table_data[56] = 16'b0101000001010000;
  assign magnitude_expected_table_data[57] = 16'b0100111110010000;
  assign magnitude_expected_table_data[58] = 16'b0101000000010000;
  assign magnitude_expected_table_data[59] = 16'b0100111111010000;
  assign magnitude_expected_table_data[60] = 16'b0100111101100000;
  assign magnitude_expected_table_data[61] = 16'b0101000001100000;
  assign magnitude_expected_table_data[62] = 16'b0100111011110000;
  assign magnitude_expected_table_data[63] = 16'b0100111111010000;
  assign magnitude_expected_table_data[64] = 16'b0100111111010000;
  assign magnitude_expected_table_data[65] = 16'b0100111011110000;
  assign magnitude_expected_table_data[66] = 16'b0101000001100000;
  assign magnitude_expected_table_data[67] = 16'b0100111101100000;
  assign magnitude_expected_table_data[68] = 16'b0100111111010000;
  assign magnitude_expected_table_data[69] = 16'b0101000000010000;
  assign magnitude_expected_table_data[70] = 16'b0100111110010000;
  assign magnitude_expected_table_data[71] = 16'b0101000001010000;
  assign magnitude_expected_table_data[72] = 16'b0101000011000000;
  assign magnitude_expected_table_data[73] = 16'b0100111100110000;
  assign magnitude_expected_table_data[74] = 16'b0101000101100000;
  assign magnitude_expected_table_data[75] = 16'b0101000100110000;
  assign magnitude_expected_table_data[76] = 16'b0100111101000000;
  assign magnitude_expected_table_data[77] = 16'b0101000100110000;
  assign magnitude_expected_table_data[78] = 16'b0101000101100000;
  assign magnitude_expected_table_data[79] = 16'b0100111100110000;
  assign magnitude_expected_table_data[80] = 16'b0101000011000000;
  assign magnitude_expected_table_data[81] = 16'b0101000001010000;
  assign magnitude_expected_table_data[82] = 16'b0100111110010000;
  assign magnitude_expected_table_data[83] = 16'b0101000000000000;
  assign magnitude_expected_table_data[84] = 16'b0100111111010000;
  assign magnitude_expected_table_data[85] = 16'b0100111101100000;
  assign magnitude_expected_table_data[86] = 16'b0101000001100000;
  assign magnitude_expected_table_data[87] = 16'b0100111011110000;
  assign magnitude_expected_table_data[88] = 16'b0100111111010000;
  assign magnitude_expected_table_data[89] = 16'b0100111111010000;
  assign magnitude_expected_table_data[90] = 16'b0100111011110000;
  assign magnitude_expected_table_data[91] = 16'b0101000001100000;
  assign magnitude_expected_table_data[92] = 16'b0100111101100000;
  assign magnitude_expected_table_data[93] = 16'b0100111111010000;
  assign magnitude_expected_table_data[94] = 16'b0101000000000000;
  assign magnitude_expected_table_data[95] = 16'b0100111110010000;
  assign magnitude_expected_table_data[96] = 16'b0101000001010000;
  assign magnitude_expected_table_data[97] = 16'b0101000011000000;
  assign magnitude_expected_table_data[98] = 16'b0100111100110000;
  assign magnitude_expected_table_data[99] = 16'b0101000101100000;
  assign magnitude_expected_table_data[100] = 16'b0101000100110000;
  assign magnitude_expected_table_data[101] = 16'b0100111101000000;
  assign magnitude_expected_table_data[102] = 16'b0101000100110000;
  assign magnitude_expected_table_data[103] = 16'b0101000101100000;
  assign magnitude_expected_table_data[104] = 16'b0100111100110000;
  assign magnitude_expected_table_data[105] = 16'b0101000011000000;
  assign magnitude_expected_table_data[106] = 16'b0101000001010000;
  assign magnitude_expected_table_data[107] = 16'b0100111110010000;
  assign magnitude_expected_table_data[108] = 16'b0101000000010000;
  assign magnitude_expected_table_data[109] = 16'b0100111111010000;
  assign magnitude_expected_table_data[110] = 16'b0100111101100000;
  assign magnitude_expected_table_data[111] = 16'b0101000001100000;
  assign magnitude_expected_table_data[112] = 16'b0100111011110000;
  assign magnitude_expected_table_data[113] = 16'b0100111111010000;
  assign magnitude_expected_table_data[114] = 16'b0100111111010000;
  assign magnitude_expected_table_data[115] = 16'b0100111011110000;
  assign magnitude_expected_table_data[116] = 16'b0101000001100000;
  assign magnitude_expected_table_data[117] = 16'b0100111101100000;
  assign magnitude_expected_table_data[118] = 16'b0100111111010000;
  assign magnitude_expected_table_data[119] = 16'b0101000000010000;
  assign magnitude_expected_table_data[120] = 16'b0100111110010000;
  assign magnitude_expected_table_data[121] = 16'b0101000001010000;
  assign magnitude_expected_table_data[122] = 16'b0101000011000000;
  assign magnitude_expected_table_data[123] = 16'b0100111100110000;
  assign magnitude_expected_table_data[124] = 16'b0101000101100000;
  assign magnitude_expected_table_data[125] = 16'b0101000100110000;
  assign magnitude_expected_table_data[126] = 16'b0100111101000000;
  assign magnitude_expected_table_data[127] = 16'b0101000100110000;
  assign magnitude_expected_table_data[128] = 16'b0101000101100000;
  assign magnitude_expected_table_data[129] = 16'b0100111100110000;
  assign magnitude_expected_table_data[130] = 16'b0101000011000000;
  assign magnitude_expected_table_data[131] = 16'b0101000001010000;
  assign magnitude_expected_table_data[132] = 16'b0100111110010000;
  assign magnitude_expected_table_data[133] = 16'b0101000000000000;
  assign magnitude_expected_table_data[134] = 16'b0100111111010000;
  assign magnitude_expected_table_data[135] = 16'b0100111101100000;
  assign magnitude_expected_table_data[136] = 16'b0101000001100000;
  assign magnitude_expected_table_data[137] = 16'b0100111011110000;
  assign magnitude_expected_table_data[138] = 16'b0100111111010000;
  assign magnitude_expected_table_data[139] = 16'b0100111111010000;
  assign magnitude_expected_table_data[140] = 16'b0100111011110000;
  assign magnitude_expected_table_data[141] = 16'b0101000001100000;
  assign magnitude_expected_table_data[142] = 16'b0100111101100000;
  assign magnitude_expected_table_data[143] = 16'b0100111111010000;
  assign magnitude_expected_table_data[144] = 16'b0101000000000000;
  assign magnitude_expected_table_data[145] = 16'b0100111110010000;
  assign magnitude_expected_table_data[146] = 16'b0101000001010000;
  assign magnitude_expected_table_data[147] = 16'b0101000011000000;
  assign magnitude_expected_table_data[148] = 16'b0100111100110000;
  assign magnitude_expected_table_data[149] = 16'b0101000101100000;
  assign magnitude_expected_table_data[150] = 16'b0101000100110000;
  assign magnitude_expected_table_data[151] = 16'b0100111101000000;
  assign magnitude_expected_table_data[152] = 16'b0101000100110000;
  assign magnitude_expected_table_data[153] = 16'b0101000101100000;
  assign magnitude_expected_table_data[154] = 16'b0100111100110000;
  assign magnitude_expected_table_data[155] = 16'b0101000011000000;
  assign magnitude_expected_table_data[156] = 16'b0101000001010000;
  assign magnitude_expected_table_data[157] = 16'b0100111110010000;
  assign magnitude_expected_table_data[158] = 16'b0101000000010000;
  assign magnitude_expected_table_data[159] = 16'b0100111111010000;
  assign magnitude_expected_table_data[160] = 16'b0100111101100000;
  assign magnitude_expected_table_data[161] = 16'b0101000001100000;
  assign magnitude_expected_table_data[162] = 16'b0100111011110000;
  assign magnitude_expected_table_data[163] = 16'b0100111111010000;
  assign magnitude_expected_table_data[164] = 16'b0100111111010000;
  assign magnitude_expected_table_data[165] = 16'b0100111011110000;
  assign magnitude_expected_table_data[166] = 16'b0101000001100000;
  assign magnitude_expected_table_data[167] = 16'b0100111101100000;
  assign magnitude_expected_table_data[168] = 16'b0100111111010000;
  assign magnitude_expected_table_data[169] = 16'b0101000000010000;
  assign magnitude_expected_table_data[170] = 16'b0100111110010000;
  assign magnitude_expected_table_data[171] = 16'b0101000001010000;
  assign magnitude_expected_table_data[172] = 16'b0101000011000000;
  assign magnitude_expected_table_data[173] = 16'b0100111100110000;
  assign magnitude_expected_table_data[174] = 16'b0101000101100000;
  assign magnitude_expected_table_data[175] = 16'b0101000100110000;
  assign magnitude_expected_table_data[176] = 16'b0100111101000000;
  assign magnitude_expected_table_data[177] = 16'b0101000100110000;
  assign magnitude_expected_table_data[178] = 16'b0101000101100000;
  assign magnitude_expected_table_data[179] = 16'b0100111100110000;
  assign magnitude_expected_table_data[180] = 16'b0101000011000000;
  assign magnitude_expected_table_data[181] = 16'b0101000001010000;
  assign magnitude_expected_table_data[182] = 16'b0100111110010000;
  assign magnitude_expected_table_data[183] = 16'b0101000000000000;
  assign magnitude_expected_table_data[184] = 16'b0100111111010000;
  assign magnitude_expected_table_data[185] = 16'b0100111101100000;
  assign magnitude_expected_table_data[186] = 16'b0101000001100000;
  assign magnitude_expected_table_data[187] = 16'b0100111011110000;
  assign magnitude_expected_table_data[188] = 16'b0100111111010000;
  assign magnitude_expected_table_data[189] = 16'b0100111111010000;
  assign magnitude_expected_table_data[190] = 16'b0100111011110000;
  assign magnitude_expected_table_data[191] = 16'b0101000001100000;
  assign magnitude_expected_table_data[192] = 16'b0100111101100000;
  assign magnitude_expected_table_data[193] = 16'b0100111111010000;
  assign magnitude_expected_table_data[194] = 16'b0101000000000000;
  assign magnitude_expected_table_data[195] = 16'b0100111110010000;
  assign magnitude_expected_table_data[196] = 16'b0101000001010000;
  assign magnitude_expected_table_data[197] = 16'b0101000011000000;
  assign magnitude_expected_table_data[198] = 16'b0100111100110000;
  assign magnitude_expected_table_data[199] = 16'b0101000101100000;
  assign magnitude_expected_table_data[200] = 16'b0101000100110000;
  assign magnitude_expected_table_data[201] = 16'b0100111101000000;
  assign magnitude_expected_table_data[202] = 16'b0101000100110000;
  assign magnitude_expected_table_data[203] = 16'b0101000101100000;
  assign magnitude_expected_table_data[204] = 16'b0100111100110000;
  assign magnitude_expected_table_data[205] = 16'b0101000011000000;
  assign magnitude_expected_table_data[206] = 16'b0101000001010000;
  assign magnitude_expected_table_data[207] = 16'b0100111110010000;
  assign magnitude_expected_table_data[208] = 16'b0101000000010000;
  assign magnitude_expected_table_data[209] = 16'b0100111111010000;
  assign magnitude_expected_table_data[210] = 16'b0100111101100000;
  assign magnitude_expected_table_data[211] = 16'b0101000001100000;
  assign magnitude_expected_table_data[212] = 16'b0100111011110000;
  assign magnitude_expected_table_data[213] = 16'b0100111111010000;
  assign magnitude_expected_table_data[214] = 16'b0100111111010000;
  assign magnitude_expected_table_data[215] = 16'b0100111011110000;
  assign magnitude_expected_table_data[216] = 16'b0101000001100000;
  assign magnitude_expected_table_data[217] = 16'b0100111101100000;
  assign magnitude_expected_table_data[218] = 16'b0100111111010000;
  assign magnitude_expected_table_data[219] = 16'b0101000000010000;
  assign magnitude_expected_table_data[220] = 16'b0100111110010000;
  assign magnitude_expected_table_data[221] = 16'b0101000001010000;
  assign magnitude_expected_table_data[222] = 16'b0101000011000000;
  assign magnitude_expected_table_data[223] = 16'b0100111100110000;
  assign magnitude_expected_table_data[224] = 16'b0101000101100000;
  assign magnitude_expected_table_data[225] = 16'b0101000100110000;
  assign magnitude_expected_table_data[226] = 16'b0100111101000000;
  assign magnitude_expected_table_data[227] = 16'b0101000100110000;
  assign magnitude_expected_table_data[228] = 16'b0101000101100000;
  assign magnitude_expected_table_data[229] = 16'b0100111100110000;
  assign magnitude_expected_table_data[230] = 16'b0101000011000000;
  assign magnitude_expected_table_data[231] = 16'b0101000001010000;
  assign magnitude_expected_table_data[232] = 16'b0100111110010000;
  assign magnitude_expected_table_data[233] = 16'b0101000000000000;
  assign magnitude_expected_table_data[234] = 16'b0100111111010000;
  assign magnitude_expected_table_data[235] = 16'b0100111101100000;
  assign magnitude_expected_table_data[236] = 16'b0101000001100000;
  assign magnitude_expected_table_data[237] = 16'b0100111011110000;
  assign magnitude_expected_table_data[238] = 16'b0100111111010000;
  assign magnitude_expected_table_data[239] = 16'b0100111111010000;
  assign magnitude_expected_table_data[240] = 16'b0100111011110000;
  assign magnitude_expected_table_data[241] = 16'b0101000001100000;
  assign magnitude_expected_table_data[242] = 16'b0100111101100000;
  assign magnitude_expected_table_data[243] = 16'b0100111111010000;
  assign magnitude_expected_table_data[244] = 16'b0101000000000000;
  assign magnitude_expected_table_data[245] = 16'b0100111110010000;
  assign magnitude_expected_table_data[246] = 16'b0101000001010000;
  assign magnitude_expected_table_data[247] = 16'b0101000011000000;
  assign magnitude_expected_table_data[248] = 16'b0100111100110000;
  assign magnitude_expected_table_data[249] = 16'b0101000101100000;
  assign magnitude_expected_table_data[250] = 16'b0101000100110000;
  assign magnitude_expected_table_data[251] = 16'b0100111101000000;
  assign magnitude_expected_table_data[252] = 16'b0101000100110000;
  assign magnitude_expected_table_data[253] = 16'b0101000101100000;
  assign magnitude_expected_table_data[254] = 16'b0100111100110000;
  assign magnitude_expected_table_data[255] = 16'b0101000011000000;
  assign magnitude_expected_table_data[256] = 16'b0101000001010000;
  assign magnitude_expected_table_data[257] = 16'b0100111110010000;
  assign magnitude_expected_table_data[258] = 16'b0101000000010000;
  assign magnitude_expected_table_data[259] = 16'b0100111111010000;
  assign magnitude_expected_table_data[260] = 16'b0100111101100000;
  assign magnitude_expected_table_data[261] = 16'b0101000001100000;
  assign magnitude_expected_table_data[262] = 16'b0100111011110000;
  assign magnitude_expected_table_data[263] = 16'b0100111111010000;
  assign magnitude_expected_table_data[264] = 16'b0100111111010000;
  assign magnitude_expected_table_data[265] = 16'b0100111011110000;
  assign magnitude_expected_table_data[266] = 16'b0101000001100000;
  assign magnitude_expected_table_data[267] = 16'b0100111101100000;
  assign magnitude_expected_table_data[268] = 16'b0100111111010000;
  assign magnitude_expected_table_data[269] = 16'b0101000000010000;
  assign magnitude_expected_table_data[270] = 16'b0100111110010000;
  assign magnitude_expected_table_data[271] = 16'b0101000001010000;
  assign magnitude_expected_table_data[272] = 16'b0101000011000000;
  assign magnitude_expected_table_data[273] = 16'b0100111100110000;
  assign magnitude_expected_table_data[274] = 16'b0101000101100000;
  assign magnitude_expected_table_data[275] = 16'b0101000100110000;
  assign magnitude_expected_table_data[276] = 16'b0001100111000000;
  assign magnitude_expected_table_data[277] = 16'b0001101010000000;
  assign magnitude_expected_table_data[278] = 16'b0001100100100000;
  assign magnitude_expected_table_data[279] = 16'b0001100110010000;
  assign magnitude_expected_table_data[280] = 16'b0001100111110000;
  assign magnitude_expected_table_data[281] = 16'b0001100100100000;
  assign magnitude_expected_table_data[282] = 16'b0001100100000000;
  assign magnitude_expected_table_data[283] = 16'b0001100010110000;
  assign magnitude_expected_table_data[284] = 16'b0001101001100000;
  assign magnitude_expected_table_data[285] = 16'b0001100010110000;
  assign magnitude_expected_table_data[286] = 16'b0001100110000000;
  assign magnitude_expected_table_data[287] = 16'b0001100100010000;
  assign magnitude_expected_table_data[288] = 16'b0001100100010000;
  assign magnitude_expected_table_data[289] = 16'b0001100100010000;
  assign magnitude_expected_table_data[290] = 16'b0001100100010000;
  assign magnitude_expected_table_data[291] = 16'b0001100110000000;
  assign magnitude_expected_table_data[292] = 16'b0001100010110000;
  assign magnitude_expected_table_data[293] = 16'b0001101001100000;
  assign magnitude_expected_table_data[294] = 16'b0001100010110000;
  assign magnitude_expected_table_data[295] = 16'b0001100100000000;
  assign magnitude_expected_table_data[296] = 16'b0001100100100000;
  assign magnitude_expected_table_data[297] = 16'b0001100111110000;
  assign magnitude_expected_table_data[298] = 16'b0001100110010000;
  assign magnitude_expected_table_data[299] = 16'b0001100100100000;
  assign magnitude_expected_table_data[300] = 16'b0001101010000000;
  assign magnitude_expected_table_data[301] = 16'b0001100111000000;
  assign magnitude_expected_table_data[302] = 16'b0001101010000000;
  assign magnitude_expected_table_data[303] = 16'b0001100100100000;
  assign magnitude_expected_table_data[304] = 16'b0001100110010000;
  assign magnitude_expected_table_data[305] = 16'b0001100111110000;
  assign magnitude_expected_table_data[306] = 16'b0001100100100000;
  assign magnitude_expected_table_data[307] = 16'b0001100100000000;
  assign magnitude_expected_table_data[308] = 16'b0001100010110000;
  assign magnitude_expected_table_data[309] = 16'b0001101001100000;
  assign magnitude_expected_table_data[310] = 16'b0001100010110000;
  assign magnitude_expected_table_data[311] = 16'b0001100110000000;
  assign magnitude_expected_table_data[312] = 16'b0001100100010000;
  assign magnitude_expected_table_data[313] = 16'b0001100100010000;
  assign magnitude_expected_table_data[314] = 16'b0001100100010000;
  assign magnitude_expected_table_data[315] = 16'b0001100100010000;
  assign magnitude_expected_table_data[316] = 16'b0001100110000000;
  assign magnitude_expected_table_data[317] = 16'b0001100010110000;
  assign magnitude_expected_table_data[318] = 16'b0001101001100000;
  assign magnitude_expected_table_data[319] = 16'b0001100010110000;
  assign magnitude_expected_table_data[320] = 16'b0001100100000000;
  assign magnitude_expected_table_data[321] = 16'b0001100100100000;
  assign magnitude_expected_table_data[322] = 16'b0001100111110000;
  assign magnitude_expected_table_data[323] = 16'b0001100110010000;
  assign magnitude_expected_table_data[324] = 16'b0001100100100000;
  assign magnitude_expected_table_data[325] = 16'b0001101010000000;
  assign magnitude_expected_table_data[326] = 16'b0001100111000000;
  assign magnitude_expected_table_data[327] = 16'b0001101010000000;
  assign magnitude_expected_table_data[328] = 16'b0001100100100000;
  assign magnitude_expected_table_data[329] = 16'b0001100110010000;
  assign magnitude_expected_table_data[330] = 16'b0001100111110000;
  assign magnitude_expected_table_data[331] = 16'b0001100100100000;
  assign magnitude_expected_table_data[332] = 16'b0001100100000000;
  assign magnitude_expected_table_data[333] = 16'b0001100010110000;
  assign magnitude_expected_table_data[334] = 16'b0001101001100000;
  assign magnitude_expected_table_data[335] = 16'b0001100010110000;
  assign magnitude_expected_table_data[336] = 16'b0001100110000000;
  assign magnitude_expected_table_data[337] = 16'b0001100100010000;
  assign magnitude_expected_table_data[338] = 16'b0001100100010000;
  assign magnitude_expected_table_data[339] = 16'b0001100100010000;
  assign magnitude_expected_table_data[340] = 16'b0001100100010000;
  assign magnitude_expected_table_data[341] = 16'b0001100110000000;
  assign magnitude_expected_table_data[342] = 16'b0001100010110000;
  assign magnitude_expected_table_data[343] = 16'b0001101001100000;
  assign magnitude_expected_table_data[344] = 16'b0001100010110000;
  assign magnitude_expected_table_data[345] = 16'b0001100100000000;
  assign magnitude_expected_table_data[346] = 16'b0001100100100000;
  assign magnitude_expected_table_data[347] = 16'b0001100111110000;
  assign magnitude_expected_table_data[348] = 16'b0001100110010000;
  assign magnitude_expected_table_data[349] = 16'b0001100100100000;
  assign magnitude_expected_table_data[350] = 16'b0001101010000000;
  assign magnitude_expected_table_data[351] = 16'b0001100111000000;
  assign magnitude_expected_table_data[352] = 16'b0001101010000000;
  assign magnitude_expected_table_data[353] = 16'b0001100100100000;
  assign magnitude_expected_table_data[354] = 16'b0001100110010000;
  assign magnitude_expected_table_data[355] = 16'b0001100111110000;
  assign magnitude_expected_table_data[356] = 16'b0001100100100000;
  assign magnitude_expected_table_data[357] = 16'b0001100100000000;
  assign magnitude_expected_table_data[358] = 16'b0001100010110000;
  assign magnitude_expected_table_data[359] = 16'b0001101001100000;
  assign magnitude_expected_table_data[360] = 16'b0001100010110000;
  assign magnitude_expected_table_data[361] = 16'b0001100110000000;
  assign magnitude_expected_table_data[362] = 16'b0001100100010000;
  assign magnitude_expected_table_data[363] = 16'b0001100100010000;
  assign magnitude_expected_table_data[364] = 16'b0001100100010000;
  assign magnitude_expected_table_data[365] = 16'b0001100100010000;
  assign magnitude_expected_table_data[366] = 16'b0001100110000000;
  assign magnitude_expected_table_data[367] = 16'b0001100010110000;
  assign magnitude_expected_table_data[368] = 16'b0001101001100000;
  assign magnitude_expected_table_data[369] = 16'b0001100010110000;
  assign magnitude_expected_table_data[370] = 16'b0001100100000000;
  assign magnitude_expected_table_data[371] = 16'b0001100100100000;
  assign magnitude_expected_table_data[372] = 16'b0001100111110000;
  assign magnitude_expected_table_data[373] = 16'b0001100110010000;
  assign magnitude_expected_table_data[374] = 16'b0001100100100000;
  assign magnitude_expected_table_data[375] = 16'b0001101010000000;
  assign magnitude_expected_table_data[376] = 16'b0001100111000000;
  assign magnitude_expected_table_data[377] = 16'b0001101010000000;
  assign magnitude_expected_table_data[378] = 16'b0001100100100000;
  assign magnitude_expected_table_data[379] = 16'b0001100110010000;
  assign magnitude_expected_table_data[380] = 16'b0001100111110000;
  assign magnitude_expected_table_data[381] = 16'b0001100100100000;
  assign magnitude_expected_table_data[382] = 16'b0001100100000000;
  assign magnitude_expected_table_data[383] = 16'b0001100010110000;
  assign magnitude_expected_table_data[384] = 16'b0001101001100000;
  assign magnitude_expected_table_data[385] = 16'b0001100010110000;
  assign magnitude_expected_table_data[386] = 16'b0001100110000000;
  assign magnitude_expected_table_data[387] = 16'b0001100100010000;
  assign magnitude_expected_table_data[388] = 16'b0001100100010000;
  assign magnitude_expected_table_data[389] = 16'b0001100100010000;
  assign magnitude_expected_table_data[390] = 16'b0001100100010000;
  assign magnitude_expected_table_data[391] = 16'b0001100110000000;
  assign magnitude_expected_table_data[392] = 16'b0001100010110000;
  assign magnitude_expected_table_data[393] = 16'b0001101001100000;
  assign magnitude_expected_table_data[394] = 16'b0001100010110000;
  assign magnitude_expected_table_data[395] = 16'b0001100100000000;
  assign magnitude_expected_table_data[396] = 16'b0001100100100000;
  assign magnitude_expected_table_data[397] = 16'b0001100111110000;
  assign magnitude_expected_table_data[398] = 16'b0001100110010000;
  assign magnitude_expected_table_data[399] = 16'b0001100100100000;
  assign magnitude_expected_table_data[400] = 16'b0001101010000000;
  assign magnitude_expected_table_data[401] = 16'b0001100111000000;
  assign magnitude_expected_table_data[402] = 16'b0001101010000000;
  assign magnitude_expected_table_data[403] = 16'b0001100100100000;
  assign magnitude_expected_table_data[404] = 16'b0001100110010000;
  assign magnitude_expected_table_data[405] = 16'b0001100111110000;
  assign magnitude_expected_table_data[406] = 16'b0001100100100000;
  assign magnitude_expected_table_data[407] = 16'b0001100100000000;
  assign magnitude_expected_table_data[408] = 16'b0001100010110000;
  assign magnitude_expected_table_data[409] = 16'b0001101001100000;
  assign magnitude_expected_table_data[410] = 16'b0001100010110000;
  assign magnitude_expected_table_data[411] = 16'b0001100110000000;
  assign magnitude_expected_table_data[412] = 16'b0001100100010000;
  assign magnitude_expected_table_data[413] = 16'b0001100100010000;
  assign magnitude_expected_table_data[414] = 16'b0001100100010000;
  assign magnitude_expected_table_data[415] = 16'b0001100100010000;
  assign magnitude_expected_table_data[416] = 16'b0001100110000000;
  assign magnitude_expected_table_data[417] = 16'b0001100010110000;
  assign magnitude_expected_table_data[418] = 16'b0001101001100000;
  assign magnitude_expected_table_data[419] = 16'b0001100010110000;
  assign magnitude_expected_table_data[420] = 16'b0001100100000000;
  assign magnitude_expected_table_data[421] = 16'b0001100100100000;
  assign magnitude_expected_table_data[422] = 16'b0001100111110000;
  assign magnitude_expected_table_data[423] = 16'b0001100110010000;
  assign magnitude_expected_table_data[424] = 16'b0001100100100000;
  assign magnitude_expected_table_data[425] = 16'b0001101010000000;
  assign magnitude_expected_table_data[426] = 16'b0001100111000000;
  assign magnitude_expected_table_data[427] = 16'b0001101010000000;
  assign magnitude_expected_table_data[428] = 16'b0001100100100000;
  assign magnitude_expected_table_data[429] = 16'b0001100110010000;
  assign magnitude_expected_table_data[430] = 16'b0001100111110000;
  assign magnitude_expected_table_data[431] = 16'b0001100100100000;
  assign magnitude_expected_table_data[432] = 16'b0001100100000000;
  assign magnitude_expected_table_data[433] = 16'b0001100010110000;
  assign magnitude_expected_table_data[434] = 16'b0001101001100000;
  assign magnitude_expected_table_data[435] = 16'b0001100010110000;
  assign magnitude_expected_table_data[436] = 16'b0001100110000000;
  assign magnitude_expected_table_data[437] = 16'b0001100100010000;
  assign magnitude_expected_table_data[438] = 16'b0001100100010000;
  assign magnitude_expected_table_data[439] = 16'b0001100100010000;
  assign magnitude_expected_table_data[440] = 16'b0001100100010000;
  assign magnitude_expected_table_data[441] = 16'b0001100110000000;
  assign magnitude_expected_table_data[442] = 16'b0001100010110000;
  assign magnitude_expected_table_data[443] = 16'b0001101001100000;
  assign magnitude_expected_table_data[444] = 16'b0001100010110000;
  assign magnitude_expected_table_data[445] = 16'b0001100100000000;
  assign magnitude_expected_table_data[446] = 16'b0001100100100000;
  assign magnitude_expected_table_data[447] = 16'b0001100111110000;
  assign magnitude_expected_table_data[448] = 16'b0001100110010000;
  assign magnitude_expected_table_data[449] = 16'b0001100100100000;
  assign magnitude_expected_table_data[450] = 16'b0001101010000000;
  assign magnitude_expected_table_data[451] = 16'b0001100111000000;
  assign magnitude_expected_table_data[452] = 16'b0001101010000000;
  assign magnitude_expected_table_data[453] = 16'b0001100100100000;
  assign magnitude_expected_table_data[454] = 16'b0001100110010000;
  assign magnitude_expected_table_data[455] = 16'b0001100111110000;
  assign magnitude_expected_table_data[456] = 16'b0001100100100000;
  assign magnitude_expected_table_data[457] = 16'b0001100100000000;
  assign magnitude_expected_table_data[458] = 16'b0001100010110000;
  assign magnitude_expected_table_data[459] = 16'b0001101001100000;
  assign magnitude_expected_table_data[460] = 16'b0001100010110000;
  assign magnitude_expected_table_data[461] = 16'b0001100110000000;
  assign magnitude_expected_table_data[462] = 16'b0001100100010000;
  assign magnitude_expected_table_data[463] = 16'b0001100100010000;
  assign magnitude_expected_table_data[464] = 16'b0001100100010000;
  assign magnitude_expected_table_data[465] = 16'b0001100100010000;
  assign magnitude_expected_table_data[466] = 16'b0001100110000000;
  assign magnitude_expected_table_data[467] = 16'b0001100010110000;
  assign magnitude_expected_table_data[468] = 16'b0001101001100000;
  assign magnitude_expected_table_data[469] = 16'b0001100010110000;
  assign magnitude_expected_table_data[470] = 16'b0001100100000000;
  assign magnitude_expected_table_data[471] = 16'b0001100100100000;
  assign magnitude_expected_table_data[472] = 16'b0001100111110000;
  assign magnitude_expected_table_data[473] = 16'b0001100110010000;
  assign magnitude_expected_table_data[474] = 16'b0001100100100000;
  assign magnitude_expected_table_data[475] = 16'b0001101010000000;
  assign magnitude_expected_table_data[476] = 16'b0001100111000000;
  assign magnitude_expected_table_data[477] = 16'b0001101010000000;
  assign magnitude_expected_table_data[478] = 16'b0001100100100000;
  assign magnitude_expected_table_data[479] = 16'b0001100110010000;
  assign magnitude_expected_table_data[480] = 16'b0001100111110000;
  assign magnitude_expected_table_data[481] = 16'b0001100100100000;
  assign magnitude_expected_table_data[482] = 16'b0001100100000000;
  assign magnitude_expected_table_data[483] = 16'b0001100010110000;
  assign magnitude_expected_table_data[484] = 16'b0001101001100000;
  assign magnitude_expected_table_data[485] = 16'b0001100010110000;
  assign magnitude_expected_table_data[486] = 16'b0001100110000000;
  assign magnitude_expected_table_data[487] = 16'b0001100100010000;
  assign magnitude_expected_table_data[488] = 16'b0001100100010000;
  assign magnitude_expected_table_data[489] = 16'b0001100100010000;
  assign magnitude_expected_table_data[490] = 16'b0001100100010000;
  assign magnitude_expected_table_data[491] = 16'b0001100110000000;
  assign magnitude_expected_table_data[492] = 16'b0001100010110000;
  assign magnitude_expected_table_data[493] = 16'b0001101001100000;
  assign magnitude_expected_table_data[494] = 16'b0001100010110000;
  assign magnitude_expected_table_data[495] = 16'b0001100100000000;
  assign magnitude_expected_table_data[496] = 16'b0001100100100000;
  assign magnitude_expected_table_data[497] = 16'b0001100111110000;
  assign magnitude_expected_table_data[498] = 16'b0001100110010000;
  assign magnitude_expected_table_data[499] = 16'b0001100100100000;
  assign magnitude_expected_table_data[500] = 16'b0001101010000000;
  assign magnitude_expected_table_data[501] = 16'b0001100111000000;
  assign magnitude_expected_table_data[502] = 16'b0001101010000000;
  assign magnitude_expected_table_data[503] = 16'b0001100100100000;
  assign magnitude_expected_table_data[504] = 16'b0001100110010000;
  assign magnitude_expected_table_data[505] = 16'b0001100111110000;
  assign magnitude_expected_table_data[506] = 16'b0001100100100000;
  assign magnitude_expected_table_data[507] = 16'b0001100100000000;
  assign magnitude_expected_table_data[508] = 16'b0001100010110000;
  assign magnitude_expected_table_data[509] = 16'b0001101001100000;
  assign magnitude_expected_table_data[510] = 16'b0001100010110000;
  assign magnitude_expected_table_data[511] = 16'b0001100110000000;
  assign magnitude_expected_table_data[512] = 16'b0001100100010000;
  assign magnitude_expected_table_data[513] = 16'b0001100100010000;
  assign magnitude_expected_table_data[514] = 16'b0001100100010000;
  assign magnitude_expected_table_data[515] = 16'b0001100100010000;
  assign magnitude_expected_table_data[516] = 16'b0001100110000000;
  assign magnitude_expected_table_data[517] = 16'b0001100010110000;
  assign magnitude_expected_table_data[518] = 16'b0001101001100000;
  assign magnitude_expected_table_data[519] = 16'b0001100010110000;
  assign magnitude_expected_table_data[520] = 16'b0001100100000000;
  assign magnitude_expected_table_data[521] = 16'b0001100100100000;
  assign magnitude_expected_table_data[522] = 16'b0001100111110000;
  assign magnitude_expected_table_data[523] = 16'b0001100110010000;
  assign magnitude_expected_table_data[524] = 16'b0001100100100000;
  assign magnitude_expected_table_data[525] = 16'b0001101010000000;
  assign magnitude_expected_table_data[526] = 16'b0010010000100000;
  assign magnitude_expected_table_data[527] = 16'b0010010010110000;
  assign magnitude_expected_table_data[528] = 16'b0010010000000000;
  assign magnitude_expected_table_data[529] = 16'b0010001110000000;
  assign magnitude_expected_table_data[530] = 16'b0010001101100000;
  assign magnitude_expected_table_data[531] = 16'b0010001100110000;
  assign magnitude_expected_table_data[532] = 16'b0010001111100000;
  assign magnitude_expected_table_data[533] = 16'b0010010011110000;
  assign magnitude_expected_table_data[534] = 16'b0010001111100000;
  assign magnitude_expected_table_data[535] = 16'b0010010000100000;
  assign magnitude_expected_table_data[536] = 16'b0010010100100000;
  assign magnitude_expected_table_data[537] = 16'b0010010000100000;
  assign magnitude_expected_table_data[538] = 16'b0010001111110000;
  assign magnitude_expected_table_data[539] = 16'b0010010000110000;
  assign magnitude_expected_table_data[540] = 16'b0010010011100000;
  assign magnitude_expected_table_data[541] = 16'b0010010011010000;
  assign magnitude_expected_table_data[542] = 16'b0010010001100000;
  assign magnitude_expected_table_data[543] = 16'b0010001111110000;
  assign magnitude_expected_table_data[544] = 16'b0010001101100000;
  assign magnitude_expected_table_data[545] = 16'b0010001111110000;
  assign magnitude_expected_table_data[546] = 16'b0010001110100000;
  assign magnitude_expected_table_data[547] = 16'b0010010000100000;
  assign magnitude_expected_table_data[548] = 16'b0010010100000000;
  assign magnitude_expected_table_data[549] = 16'b0010001111100000;
  assign magnitude_expected_table_data[550] = 16'b0010001110110000;
  assign magnitude_expected_table_data[551] = 16'b0010010000100000;
  assign magnitude_expected_table_data[552] = 16'b0010010010110000;
  assign magnitude_expected_table_data[553] = 16'b0010010000000000;
  assign magnitude_expected_table_data[554] = 16'b0010001110000000;
  assign magnitude_expected_table_data[555] = 16'b0010001101100000;
  assign magnitude_expected_table_data[556] = 16'b0010001100110000;
  assign magnitude_expected_table_data[557] = 16'b0010001111100000;
  assign magnitude_expected_table_data[558] = 16'b0010010011110000;
  assign magnitude_expected_table_data[559] = 16'b0010001111100000;
  assign magnitude_expected_table_data[560] = 16'b0010010000100000;
  assign magnitude_expected_table_data[561] = 16'b0010010100100000;
  assign magnitude_expected_table_data[562] = 16'b0010010000100000;
  assign magnitude_expected_table_data[563] = 16'b0010001111110000;
  assign magnitude_expected_table_data[564] = 16'b0010010000110000;
  assign magnitude_expected_table_data[565] = 16'b0010010011100000;
  assign magnitude_expected_table_data[566] = 16'b0010010011010000;
  assign magnitude_expected_table_data[567] = 16'b0010010001100000;
  assign magnitude_expected_table_data[568] = 16'b0010001111110000;
  assign magnitude_expected_table_data[569] = 16'b0010001101100000;
  assign magnitude_expected_table_data[570] = 16'b0010001111110000;
  assign magnitude_expected_table_data[571] = 16'b0010001110100000;
  assign magnitude_expected_table_data[572] = 16'b0010010000100000;
  assign magnitude_expected_table_data[573] = 16'b0010010100000000;
  assign magnitude_expected_table_data[574] = 16'b0010001111100000;
  assign magnitude_expected_table_data[575] = 16'b0010001110110000;
  assign magnitude_expected_table_data[576] = 16'b0010010000100000;
  assign magnitude_expected_table_data[577] = 16'b0010010010110000;
  assign magnitude_expected_table_data[578] = 16'b0010010000000000;
  assign magnitude_expected_table_data[579] = 16'b0010001110000000;
  assign magnitude_expected_table_data[580] = 16'b0010001101100000;
  assign magnitude_expected_table_data[581] = 16'b0010001100110000;
  assign magnitude_expected_table_data[582] = 16'b0010001111100000;
  assign magnitude_expected_table_data[583] = 16'b0010010011110000;
  assign magnitude_expected_table_data[584] = 16'b0010001111100000;
  assign magnitude_expected_table_data[585] = 16'b0010010000100000;
  assign magnitude_expected_table_data[586] = 16'b0010010100100000;
  assign magnitude_expected_table_data[587] = 16'b0010010000100000;
  assign magnitude_expected_table_data[588] = 16'b0010001111110000;
  assign magnitude_expected_table_data[589] = 16'b0010010000110000;
  assign magnitude_expected_table_data[590] = 16'b0010010011100000;
  assign magnitude_expected_table_data[591] = 16'b0010010011010000;
  assign magnitude_expected_table_data[592] = 16'b0010010001100000;
  assign magnitude_expected_table_data[593] = 16'b0010001111110000;
  assign magnitude_expected_table_data[594] = 16'b0010001101100000;
  assign magnitude_expected_table_data[595] = 16'b0010001111110000;
  assign magnitude_expected_table_data[596] = 16'b0010001110100000;
  assign magnitude_expected_table_data[597] = 16'b0010010000100000;
  assign magnitude_expected_table_data[598] = 16'b0010010100000000;
  assign magnitude_expected_table_data[599] = 16'b0010001111100000;
  assign magnitude_expected_table_data[600] = 16'b0010001110110000;
  assign magnitude_expected_table_data[601] = 16'b0010010000100000;
  assign magnitude_expected_table_data[602] = 16'b0010010010110000;
  assign magnitude_expected_table_data[603] = 16'b0010010000000000;
  assign magnitude_expected_table_data[604] = 16'b0010001110000000;
  assign magnitude_expected_table_data[605] = 16'b0010001101100000;
  assign magnitude_expected_table_data[606] = 16'b0010001100110000;
  assign magnitude_expected_table_data[607] = 16'b0010001111100000;
  assign magnitude_expected_table_data[608] = 16'b0010010011110000;
  assign magnitude_expected_table_data[609] = 16'b0010001111100000;
  assign magnitude_expected_table_data[610] = 16'b0010010000100000;
  assign magnitude_expected_table_data[611] = 16'b0010010100100000;
  assign magnitude_expected_table_data[612] = 16'b0010010000100000;
  assign magnitude_expected_table_data[613] = 16'b0010001111110000;
  assign magnitude_expected_table_data[614] = 16'b0010010000110000;
  assign magnitude_expected_table_data[615] = 16'b0010010011100000;
  assign magnitude_expected_table_data[616] = 16'b0010010011010000;
  assign magnitude_expected_table_data[617] = 16'b0010010001100000;
  assign magnitude_expected_table_data[618] = 16'b0010001111110000;
  assign magnitude_expected_table_data[619] = 16'b0010001101100000;
  assign magnitude_expected_table_data[620] = 16'b0010001111110000;
  assign magnitude_expected_table_data[621] = 16'b0010001110100000;
  assign magnitude_expected_table_data[622] = 16'b0010010000100000;
  assign magnitude_expected_table_data[623] = 16'b0010010100000000;
  assign magnitude_expected_table_data[624] = 16'b0010001111100000;
  assign magnitude_expected_table_data[625] = 16'b0010001110110000;
  assign magnitude_expected_table_data[626] = 16'b0010010000100000;
  assign magnitude_expected_table_data[627] = 16'b0010010010110000;
  assign magnitude_expected_table_data[628] = 16'b0010010000000000;
  assign magnitude_expected_table_data[629] = 16'b0010001110000000;
  assign magnitude_expected_table_data[630] = 16'b0010001101100000;
  assign magnitude_expected_table_data[631] = 16'b0010001100110000;
  assign magnitude_expected_table_data[632] = 16'b0010001111100000;
  assign magnitude_expected_table_data[633] = 16'b0010010011110000;
  assign magnitude_expected_table_data[634] = 16'b0010001111100000;
  assign magnitude_expected_table_data[635] = 16'b0010010000100000;
  assign magnitude_expected_table_data[636] = 16'b0010010100100000;
  assign magnitude_expected_table_data[637] = 16'b0010010000100000;
  assign magnitude_expected_table_data[638] = 16'b0010001111110000;
  assign magnitude_expected_table_data[639] = 16'b0010010000110000;
  assign magnitude_expected_table_data[640] = 16'b0010010011100000;
  assign magnitude_expected_table_data[641] = 16'b0010010011010000;
  assign magnitude_expected_table_data[642] = 16'b0010010001100000;
  assign magnitude_expected_table_data[643] = 16'b0010001111110000;
  assign magnitude_expected_table_data[644] = 16'b0010001101100000;
  assign magnitude_expected_table_data[645] = 16'b0010001111110000;
  assign magnitude_expected_table_data[646] = 16'b0010001110100000;
  assign magnitude_expected_table_data[647] = 16'b0010010000100000;
  assign magnitude_expected_table_data[648] = 16'b0010010100000000;
  assign magnitude_expected_table_data[649] = 16'b0010001111100000;
  assign magnitude_expected_table_data[650] = 16'b0010001110110000;
  assign magnitude_expected_table_data[651] = 16'b0010010000100000;
  assign magnitude_expected_table_data[652] = 16'b0010010010110000;
  assign magnitude_expected_table_data[653] = 16'b0010010000000000;
  assign magnitude_expected_table_data[654] = 16'b0010001110000000;
  assign magnitude_expected_table_data[655] = 16'b0010001101100000;
  assign magnitude_expected_table_data[656] = 16'b0010001100110000;
  assign magnitude_expected_table_data[657] = 16'b0010001111100000;
  assign magnitude_expected_table_data[658] = 16'b0010010011110000;
  assign magnitude_expected_table_data[659] = 16'b0010001111100000;
  assign magnitude_expected_table_data[660] = 16'b0010010000100000;
  assign magnitude_expected_table_data[661] = 16'b0010010100100000;
  assign magnitude_expected_table_data[662] = 16'b0010010000100000;
  assign magnitude_expected_table_data[663] = 16'b0010001111110000;
  assign magnitude_expected_table_data[664] = 16'b0010010000110000;
  assign magnitude_expected_table_data[665] = 16'b0010010011100000;
  assign magnitude_expected_table_data[666] = 16'b0010010011010000;
  assign magnitude_expected_table_data[667] = 16'b0010010001100000;
  assign magnitude_expected_table_data[668] = 16'b0010001111110000;
  assign magnitude_expected_table_data[669] = 16'b0010001101100000;
  assign magnitude_expected_table_data[670] = 16'b0010001111110000;
  assign magnitude_expected_table_data[671] = 16'b0010001110100000;
  assign magnitude_expected_table_data[672] = 16'b0010010000100000;
  assign magnitude_expected_table_data[673] = 16'b0010010100000000;
  assign magnitude_expected_table_data[674] = 16'b0010001111100000;
  assign magnitude_expected_table_data[675] = 16'b0010001110110000;
  assign magnitude_expected_table_data[676] = 16'b0010010000100000;
  assign magnitude_expected_table_data[677] = 16'b0010010010110000;
  assign magnitude_expected_table_data[678] = 16'b0010010000000000;
  assign magnitude_expected_table_data[679] = 16'b0010001110000000;
  assign magnitude_expected_table_data[680] = 16'b0010001101100000;
  assign magnitude_expected_table_data[681] = 16'b0010001100110000;
  assign magnitude_expected_table_data[682] = 16'b0010001111100000;
  assign magnitude_expected_table_data[683] = 16'b0010010011110000;
  assign magnitude_expected_table_data[684] = 16'b0010001111100000;
  assign magnitude_expected_table_data[685] = 16'b0010010000100000;
  assign magnitude_expected_table_data[686] = 16'b0010010100100000;
  assign magnitude_expected_table_data[687] = 16'b0010010000100000;
  assign magnitude_expected_table_data[688] = 16'b0010001111110000;
  assign magnitude_expected_table_data[689] = 16'b0010010000110000;
  assign magnitude_expected_table_data[690] = 16'b0010010011100000;
  assign magnitude_expected_table_data[691] = 16'b0010010011010000;
  assign magnitude_expected_table_data[692] = 16'b0010010001100000;
  assign magnitude_expected_table_data[693] = 16'b0010001111110000;
  assign magnitude_expected_table_data[694] = 16'b0010001101100000;
  assign magnitude_expected_table_data[695] = 16'b0010001111110000;
  assign magnitude_expected_table_data[696] = 16'b0010001110100000;
  assign magnitude_expected_table_data[697] = 16'b0010010000100000;
  assign magnitude_expected_table_data[698] = 16'b0010010100000000;
  assign magnitude_expected_table_data[699] = 16'b0010001111100000;
  assign magnitude_expected_table_data[700] = 16'b0010001110110000;
  assign magnitude_expected_table_data[701] = 16'b0010010000100000;
  assign magnitude_expected_table_data[702] = 16'b0010010010110000;
  assign magnitude_expected_table_data[703] = 16'b0010010000000000;
  assign magnitude_expected_table_data[704] = 16'b0010001110000000;
  assign magnitude_expected_table_data[705] = 16'b0010001101100000;
  assign magnitude_expected_table_data[706] = 16'b0010001100110000;
  assign magnitude_expected_table_data[707] = 16'b0010001111100000;
  assign magnitude_expected_table_data[708] = 16'b0010010011110000;
  assign magnitude_expected_table_data[709] = 16'b0010001111100000;
  assign magnitude_expected_table_data[710] = 16'b0010010000100000;
  assign magnitude_expected_table_data[711] = 16'b0010010100100000;
  assign magnitude_expected_table_data[712] = 16'b0010010000100000;
  assign magnitude_expected_table_data[713] = 16'b0010001111110000;
  assign magnitude_expected_table_data[714] = 16'b0010010000110000;
  assign magnitude_expected_table_data[715] = 16'b0010010011100000;
  assign magnitude_expected_table_data[716] = 16'b0010010011010000;
  assign magnitude_expected_table_data[717] = 16'b0010010001100000;
  assign magnitude_expected_table_data[718] = 16'b0010001111110000;
  assign magnitude_expected_table_data[719] = 16'b0010001101100000;
  assign magnitude_expected_table_data[720] = 16'b0010001111110000;
  assign magnitude_expected_table_data[721] = 16'b0010001110100000;
  assign magnitude_expected_table_data[722] = 16'b0010010000100000;
  assign magnitude_expected_table_data[723] = 16'b0010010100000000;
  assign magnitude_expected_table_data[724] = 16'b0010001111100000;
  assign magnitude_expected_table_data[725] = 16'b0010001110110000;
  assign magnitude_expected_table_data[726] = 16'b0010010000100000;
  assign magnitude_expected_table_data[727] = 16'b0010010010110000;
  assign magnitude_expected_table_data[728] = 16'b0010010000000000;
  assign magnitude_expected_table_data[729] = 16'b0010001110000000;
  assign magnitude_expected_table_data[730] = 16'b0010001101100000;
  assign magnitude_expected_table_data[731] = 16'b0010001100110000;
  assign magnitude_expected_table_data[732] = 16'b0010001111100000;
  assign magnitude_expected_table_data[733] = 16'b0010010011110000;
  assign magnitude_expected_table_data[734] = 16'b0010001111100000;
  assign magnitude_expected_table_data[735] = 16'b0010010000100000;
  assign magnitude_expected_table_data[736] = 16'b0010010100100000;
  assign magnitude_expected_table_data[737] = 16'b0010010000100000;
  assign magnitude_expected_table_data[738] = 16'b0010001111110000;
  assign magnitude_expected_table_data[739] = 16'b0010010000110000;
  assign magnitude_expected_table_data[740] = 16'b0010010011100000;
  assign magnitude_expected_table_data[741] = 16'b0010010011010000;
  assign magnitude_expected_table_data[742] = 16'b0010010001100000;
  assign magnitude_expected_table_data[743] = 16'b0010001111110000;
  assign magnitude_expected_table_data[744] = 16'b0010001101100000;
  assign magnitude_expected_table_data[745] = 16'b0010001111110000;
  assign magnitude_expected_table_data[746] = 16'b0010001110100000;
  assign magnitude_expected_table_data[747] = 16'b0010010000100000;
  assign magnitude_expected_table_data[748] = 16'b0010010100000000;
  assign magnitude_expected_table_data[749] = 16'b0010001111100000;
  assign magnitude_expected_table_data[750] = 16'b0010001110110000;
  assign magnitude_expected_table_data[751] = 16'b0010010000100000;
  assign magnitude_expected_table_data[752] = 16'b0010010010110000;
  assign magnitude_expected_table_data[753] = 16'b0010010000000000;
  assign magnitude_expected_table_data[754] = 16'b0010001110000000;
  assign magnitude_expected_table_data[755] = 16'b0010001101100000;
  assign magnitude_expected_table_data[756] = 16'b0010001100110000;
  assign magnitude_expected_table_data[757] = 16'b0010001111100000;
  assign magnitude_expected_table_data[758] = 16'b0010010011110000;
  assign magnitude_expected_table_data[759] = 16'b0010001111100000;
  assign magnitude_expected_table_data[760] = 16'b0010010000100000;
  assign magnitude_expected_table_data[761] = 16'b0010010100100000;
  assign magnitude_expected_table_data[762] = 16'b0010010000100000;
  assign magnitude_expected_table_data[763] = 16'b0010001111110000;
  assign magnitude_expected_table_data[764] = 16'b0010010000110000;
  assign magnitude_expected_table_data[765] = 16'b0010010011100000;
  assign magnitude_expected_table_data[766] = 16'b0010010011010000;
  assign magnitude_expected_table_data[767] = 16'b0010010001100000;
  assign magnitude_expected_table_data[768] = 16'b0010001111110000;
  assign magnitude_expected_table_data[769] = 16'b0010001101100000;
  assign magnitude_expected_table_data[770] = 16'b0010001111110000;
  assign magnitude_expected_table_data[771] = 16'b0010001110100000;
  assign magnitude_expected_table_data[772] = 16'b0010010000100000;
  assign magnitude_expected_table_data[773] = 16'b0010010100000000;
  assign magnitude_expected_table_data[774] = 16'b0010001111100000;
  assign magnitude_expected_table_data[775] = 16'b0010001110110000;
  assign magnitude_expected_table_data[776] = 16'b0000001101100000;
  assign magnitude_expected_table_data[777] = 16'b0000001010010000;
  assign magnitude_expected_table_data[778] = 16'b0000001011010000;
  assign magnitude_expected_table_data[779] = 16'b0000001010110000;
  assign magnitude_expected_table_data[780] = 16'b0000001100010000;
  assign magnitude_expected_table_data[781] = 16'b0000001100010000;
  assign magnitude_expected_table_data[782] = 16'b0000010001000000;
  assign magnitude_expected_table_data[783] = 16'b0000001111000000;
  assign magnitude_expected_table_data[784] = 16'b0000001010100000;
  assign magnitude_expected_table_data[785] = 16'b0000001100000000;
  assign magnitude_expected_table_data[786] = 16'b0000001010010000;
  assign magnitude_expected_table_data[787] = 16'b0000001111010000;
  assign magnitude_expected_table_data[788] = 16'b0000010000100000;
  assign magnitude_expected_table_data[789] = 16'b0000001100100000;
  assign magnitude_expected_table_data[790] = 16'b0000001011110000;
  assign magnitude_expected_table_data[791] = 16'b0000001011000000;
  assign magnitude_expected_table_data[792] = 16'b0000001010010000;
  assign magnitude_expected_table_data[793] = 16'b0000001010100000;
  assign magnitude_expected_table_data[794] = 16'b0000001001110000;
  assign magnitude_expected_table_data[795] = 16'b0000001100100000;
  assign magnitude_expected_table_data[796] = 16'b0000010010000000;
  assign magnitude_expected_table_data[797] = 16'b0000010000010000;
  assign magnitude_expected_table_data[798] = 16'b0000001111110000;
  assign magnitude_expected_table_data[799] = 16'b0000010000010000;
  assign magnitude_expected_table_data[800] = 16'b0000010010010000;
  assign magnitude_expected_table_data[801] = 16'b0000001101100000;
  assign magnitude_expected_table_data[802] = 16'b0000001010010000;
  assign magnitude_expected_table_data[803] = 16'b0000001011010000;
  assign magnitude_expected_table_data[804] = 16'b0000001010110000;
  assign magnitude_expected_table_data[805] = 16'b0000001100010000;
  assign magnitude_expected_table_data[806] = 16'b0000001100010000;
  assign magnitude_expected_table_data[807] = 16'b0000010001000000;
  assign magnitude_expected_table_data[808] = 16'b0000001111000000;
  assign magnitude_expected_table_data[809] = 16'b0000001010100000;
  assign magnitude_expected_table_data[810] = 16'b0000001100000000;
  assign magnitude_expected_table_data[811] = 16'b0000001010010000;
  assign magnitude_expected_table_data[812] = 16'b0000001111010000;
  assign magnitude_expected_table_data[813] = 16'b0000010000100000;
  assign magnitude_expected_table_data[814] = 16'b0000001100100000;
  assign magnitude_expected_table_data[815] = 16'b0000001011110000;
  assign magnitude_expected_table_data[816] = 16'b0000001011000000;
  assign magnitude_expected_table_data[817] = 16'b0000001010010000;
  assign magnitude_expected_table_data[818] = 16'b0000001010100000;
  assign magnitude_expected_table_data[819] = 16'b0000001001110000;
  assign magnitude_expected_table_data[820] = 16'b0000001100100000;
  assign magnitude_expected_table_data[821] = 16'b0000010010000000;
  assign magnitude_expected_table_data[822] = 16'b0000010000010000;
  assign magnitude_expected_table_data[823] = 16'b0000001111110000;
  assign magnitude_expected_table_data[824] = 16'b0000010000010000;
  assign magnitude_expected_table_data[825] = 16'b0000010010010000;
  assign magnitude_expected_table_data[826] = 16'b0000001101100000;
  assign magnitude_expected_table_data[827] = 16'b0000001010010000;
  assign magnitude_expected_table_data[828] = 16'b0000001011010000;
  assign magnitude_expected_table_data[829] = 16'b0000001010110000;
  assign magnitude_expected_table_data[830] = 16'b0000001100010000;
  assign magnitude_expected_table_data[831] = 16'b0000001100010000;
  assign magnitude_expected_table_data[832] = 16'b0000010001000000;
  assign magnitude_expected_table_data[833] = 16'b0000001111000000;
  assign magnitude_expected_table_data[834] = 16'b0000001010100000;
  assign magnitude_expected_table_data[835] = 16'b0000001100000000;
  assign magnitude_expected_table_data[836] = 16'b0000001010010000;
  assign magnitude_expected_table_data[837] = 16'b0000001111010000;
  assign magnitude_expected_table_data[838] = 16'b0000010000100000;
  assign magnitude_expected_table_data[839] = 16'b0000001100100000;
  assign magnitude_expected_table_data[840] = 16'b0000001011110000;
  assign magnitude_expected_table_data[841] = 16'b0000001011000000;
  assign magnitude_expected_table_data[842] = 16'b0000001010010000;
  assign magnitude_expected_table_data[843] = 16'b0000001010100000;
  assign magnitude_expected_table_data[844] = 16'b0000001001110000;
  assign magnitude_expected_table_data[845] = 16'b0000001100100000;
  assign magnitude_expected_table_data[846] = 16'b0000010010000000;
  assign magnitude_expected_table_data[847] = 16'b0000010000010000;
  assign magnitude_expected_table_data[848] = 16'b0000001111110000;
  assign magnitude_expected_table_data[849] = 16'b0000010000010000;
  assign magnitude_expected_table_data[850] = 16'b0000010010010000;
  assign magnitude_expected_table_data[851] = 16'b0000001101100000;
  assign magnitude_expected_table_data[852] = 16'b0000001010010000;
  assign magnitude_expected_table_data[853] = 16'b0000001011010000;
  assign magnitude_expected_table_data[854] = 16'b0000001010110000;
  assign magnitude_expected_table_data[855] = 16'b0000001100010000;
  assign magnitude_expected_table_data[856] = 16'b0000001100010000;
  assign magnitude_expected_table_data[857] = 16'b0000010001000000;
  assign magnitude_expected_table_data[858] = 16'b0000001111000000;
  assign magnitude_expected_table_data[859] = 16'b0000001010100000;
  assign magnitude_expected_table_data[860] = 16'b0000001100000000;
  assign magnitude_expected_table_data[861] = 16'b0000001010010000;
  assign magnitude_expected_table_data[862] = 16'b0000001111010000;
  assign magnitude_expected_table_data[863] = 16'b0000010000100000;
  assign magnitude_expected_table_data[864] = 16'b0000001100100000;
  assign magnitude_expected_table_data[865] = 16'b0000001011110000;
  assign magnitude_expected_table_data[866] = 16'b0000001011000000;
  assign magnitude_expected_table_data[867] = 16'b0000001010010000;
  assign magnitude_expected_table_data[868] = 16'b0000001010100000;
  assign magnitude_expected_table_data[869] = 16'b0000001001110000;
  assign magnitude_expected_table_data[870] = 16'b0000001100100000;
  assign magnitude_expected_table_data[871] = 16'b0000010010000000;
  assign magnitude_expected_table_data[872] = 16'b0000010000010000;
  assign magnitude_expected_table_data[873] = 16'b0000001111110000;
  assign magnitude_expected_table_data[874] = 16'b0000010000010000;
  assign magnitude_expected_table_data[875] = 16'b0000010010010000;
  assign magnitude_expected_table_data[876] = 16'b0000001101100000;
  assign magnitude_expected_table_data[877] = 16'b0000001010010000;
  assign magnitude_expected_table_data[878] = 16'b0000001011010000;
  assign magnitude_expected_table_data[879] = 16'b0000001010110000;
  assign magnitude_expected_table_data[880] = 16'b0000001100010000;
  assign magnitude_expected_table_data[881] = 16'b0000001100010000;
  assign magnitude_expected_table_data[882] = 16'b0000010001000000;
  assign magnitude_expected_table_data[883] = 16'b0000001111000000;
  assign magnitude_expected_table_data[884] = 16'b0000001010100000;
  assign magnitude_expected_table_data[885] = 16'b0000001100000000;
  assign magnitude_expected_table_data[886] = 16'b0000001010010000;
  assign magnitude_expected_table_data[887] = 16'b0000001111010000;
  assign magnitude_expected_table_data[888] = 16'b0000010000100000;
  assign magnitude_expected_table_data[889] = 16'b0000001100100000;
  assign magnitude_expected_table_data[890] = 16'b0000001011110000;
  assign magnitude_expected_table_data[891] = 16'b0000001011000000;
  assign magnitude_expected_table_data[892] = 16'b0000001010010000;
  assign magnitude_expected_table_data[893] = 16'b0000001010100000;
  assign magnitude_expected_table_data[894] = 16'b0000001001110000;
  assign magnitude_expected_table_data[895] = 16'b0000001100100000;
  assign magnitude_expected_table_data[896] = 16'b0000010010000000;
  assign magnitude_expected_table_data[897] = 16'b0000010000010000;
  assign magnitude_expected_table_data[898] = 16'b0000001111110000;
  assign magnitude_expected_table_data[899] = 16'b0000010000010000;
  assign magnitude_expected_table_data[900] = 16'b0000010010010000;
  assign magnitude_expected_table_data[901] = 16'b0000001101100000;
  assign magnitude_expected_table_data[902] = 16'b0000001010010000;
  assign magnitude_expected_table_data[903] = 16'b0000001011010000;
  assign magnitude_expected_table_data[904] = 16'b0000001010110000;
  assign magnitude_expected_table_data[905] = 16'b0000001100010000;
  assign magnitude_expected_table_data[906] = 16'b0000001100010000;
  assign magnitude_expected_table_data[907] = 16'b0000010001000000;
  assign magnitude_expected_table_data[908] = 16'b0000001111000000;
  assign magnitude_expected_table_data[909] = 16'b0000001010100000;
  assign magnitude_expected_table_data[910] = 16'b0000001100000000;
  assign magnitude_expected_table_data[911] = 16'b0000001010010000;
  assign magnitude_expected_table_data[912] = 16'b0000001111010000;
  assign magnitude_expected_table_data[913] = 16'b0000010000100000;
  assign magnitude_expected_table_data[914] = 16'b0000001100100000;
  assign magnitude_expected_table_data[915] = 16'b0000001011110000;
  assign magnitude_expected_table_data[916] = 16'b0000001011000000;
  assign magnitude_expected_table_data[917] = 16'b0000001010010000;
  assign magnitude_expected_table_data[918] = 16'b0000001010100000;
  assign magnitude_expected_table_data[919] = 16'b0000001001110000;
  assign magnitude_expected_table_data[920] = 16'b0000001100100000;
  assign magnitude_expected_table_data[921] = 16'b0000010010000000;
  assign magnitude_expected_table_data[922] = 16'b0000010000010000;
  assign magnitude_expected_table_data[923] = 16'b0000001111110000;
  assign magnitude_expected_table_data[924] = 16'b0000010000010000;
  assign magnitude_expected_table_data[925] = 16'b0000010010010000;
  assign magnitude_expected_table_data[926] = 16'b0000001101100000;
  assign magnitude_expected_table_data[927] = 16'b0000001010010000;
  assign magnitude_expected_table_data[928] = 16'b0000001011010000;
  assign magnitude_expected_table_data[929] = 16'b0000001010110000;
  assign magnitude_expected_table_data[930] = 16'b0000001100010000;
  assign magnitude_expected_table_data[931] = 16'b0000001100010000;
  assign magnitude_expected_table_data[932] = 16'b0000010001000000;
  assign magnitude_expected_table_data[933] = 16'b0000001111000000;
  assign magnitude_expected_table_data[934] = 16'b0000001010100000;
  assign magnitude_expected_table_data[935] = 16'b0000001100000000;
  assign magnitude_expected_table_data[936] = 16'b0000001010010000;
  assign magnitude_expected_table_data[937] = 16'b0000001111010000;
  assign magnitude_expected_table_data[938] = 16'b0000010000100000;
  assign magnitude_expected_table_data[939] = 16'b0000001100100000;
  assign magnitude_expected_table_data[940] = 16'b0000001011110000;
  assign magnitude_expected_table_data[941] = 16'b0000001011000000;
  assign magnitude_expected_table_data[942] = 16'b0000001010010000;
  assign magnitude_expected_table_data[943] = 16'b0000001010100000;
  assign magnitude_expected_table_data[944] = 16'b0000001001110000;
  assign magnitude_expected_table_data[945] = 16'b0000001100100000;
  assign magnitude_expected_table_data[946] = 16'b0000010010000000;
  assign magnitude_expected_table_data[947] = 16'b0000010000010000;
  assign magnitude_expected_table_data[948] = 16'b0000001111110000;
  assign magnitude_expected_table_data[949] = 16'b0000010000010000;
  assign magnitude_expected_table_data[950] = 16'b0000010010010000;
  assign magnitude_expected_table_data[951] = 16'b0000001101100000;
  assign magnitude_expected_table_data[952] = 16'b0000001010010000;
  assign magnitude_expected_table_data[953] = 16'b0000001011010000;
  assign magnitude_expected_table_data[954] = 16'b0000001010110000;
  assign magnitude_expected_table_data[955] = 16'b0000001100010000;
  assign magnitude_expected_table_data[956] = 16'b0000001100010000;
  assign magnitude_expected_table_data[957] = 16'b0000010001000000;
  assign magnitude_expected_table_data[958] = 16'b0000001111000000;
  assign magnitude_expected_table_data[959] = 16'b0000001010100000;
  assign magnitude_expected_table_data[960] = 16'b0000001100000000;
  assign magnitude_expected_table_data[961] = 16'b0000001010010000;
  assign magnitude_expected_table_data[962] = 16'b0000001111010000;
  assign magnitude_expected_table_data[963] = 16'b0000010000100000;
  assign magnitude_expected_table_data[964] = 16'b0000001100100000;
  assign magnitude_expected_table_data[965] = 16'b0000001011110000;
  assign magnitude_expected_table_data[966] = 16'b0000001011000000;
  assign magnitude_expected_table_data[967] = 16'b0000001010010000;
  assign magnitude_expected_table_data[968] = 16'b0000001010100000;
  assign magnitude_expected_table_data[969] = 16'b0000001001110000;
  assign magnitude_expected_table_data[970] = 16'b0000001100100000;
  assign magnitude_expected_table_data[971] = 16'b0000010010000000;
  assign magnitude_expected_table_data[972] = 16'b0000010000010000;
  assign magnitude_expected_table_data[973] = 16'b0000001111110000;
  assign magnitude_expected_table_data[974] = 16'b0000010000010000;
  assign magnitude_expected_table_data[975] = 16'b0000010010010000;
  assign magnitude_expected_table_data[976] = 16'b0000001101100000;
  assign magnitude_expected_table_data[977] = 16'b0000001010010000;
  assign magnitude_expected_table_data[978] = 16'b0000001011010000;
  assign magnitude_expected_table_data[979] = 16'b0000001010110000;
  assign magnitude_expected_table_data[980] = 16'b0000001100010000;
  assign magnitude_expected_table_data[981] = 16'b0000001100010000;
  assign magnitude_expected_table_data[982] = 16'b0000010001000000;
  assign magnitude_expected_table_data[983] = 16'b0000001111000000;
  assign magnitude_expected_table_data[984] = 16'b0000001010100000;
  assign magnitude_expected_table_data[985] = 16'b0000001100000000;
  assign magnitude_expected_table_data[986] = 16'b0000001010010000;
  assign magnitude_expected_table_data[987] = 16'b0000001111010000;
  assign magnitude_expected_table_data[988] = 16'b0000010000100000;
  assign magnitude_expected_table_data[989] = 16'b0000001100100000;
  assign magnitude_expected_table_data[990] = 16'b0000001011110000;
  assign magnitude_expected_table_data[991] = 16'b0000001011000000;
  assign magnitude_expected_table_data[992] = 16'b0000001010010000;
  assign magnitude_expected_table_data[993] = 16'b0000001010100000;
  assign magnitude_expected_table_data[994] = 16'b0000001001110000;
  assign magnitude_expected_table_data[995] = 16'b0000001100100000;
  assign magnitude_expected_table_data[996] = 16'b0000010010000000;
  assign magnitude_expected_table_data[997] = 16'b0000010000010000;
  assign magnitude_expected_table_data[998] = 16'b0000001111110000;
  assign magnitude_expected_table_data[999] = 16'b0000010000010000;
  assign magnitude_expected_table_data[1000] = 16'b0000010010010000;
  assign magnitude_expected_1 = magnitude_expected_table_data[magnitude_addr];



  assign magnitude_expected_2 = magnitude_expected_1;



  assign magnitude_ref = magnitude_expected_2;

  always @(posedge clk)
    begin : magnitude_checker
      if (reset_x == 1'b1) begin
        magnitude_testFailure <= 1'b0;
      end
      else begin
        if (clk_enable == 1'b1 && magnitude !== magnitude_ref) begin
          magnitude_testFailure <= 1'b1;
          $display("ERROR in magnitude at time %t : Expected '%h' Actual '%h'", $time, magnitude_ref, magnitude);
        end
      end
    end

  // Data source for alpha_arctangen_expected
  assign alpha_arctangen_expected_table_data[0] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[1] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[2] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[3] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[4] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[5] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[6] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[7] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[8] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[9] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[10] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[11] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[12] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[13] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[14] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[15] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[16] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[17] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[18] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[19] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[20] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[21] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[22] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[23] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[24] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[25] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[26] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[27] = 8'b00000100;
  assign alpha_arctangen_expected_table_data[28] = 8'b00001000;
  assign alpha_arctangen_expected_table_data[29] = 8'b00001100;
  assign alpha_arctangen_expected_table_data[30] = 8'b00010000;
  assign alpha_arctangen_expected_table_data[31] = 8'b00010101;
  assign alpha_arctangen_expected_table_data[32] = 8'b00011000;
  assign alpha_arctangen_expected_table_data[33] = 8'b00010111;
  assign alpha_arctangen_expected_table_data[34] = 8'b00010101;
  assign alpha_arctangen_expected_table_data[35] = 8'b00010100;
  assign alpha_arctangen_expected_table_data[36] = 8'b00011000;
  assign alpha_arctangen_expected_table_data[37] = 8'b00100000;
  assign alpha_arctangen_expected_table_data[38] = 8'b00101010;
  assign alpha_arctangen_expected_table_data[39] = 8'b00111011;
  assign alpha_arctangen_expected_table_data[40] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[41] = 8'b01001101;
  assign alpha_arctangen_expected_table_data[42] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[43] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[44] = 8'b01001110;
  assign alpha_arctangen_expected_table_data[45] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[46] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[47] = 8'b01010100;
  assign alpha_arctangen_expected_table_data[48] = 8'b01011000;
  assign alpha_arctangen_expected_table_data[49] = 8'b01011100;
  assign alpha_arctangen_expected_table_data[50] = 8'b01100001;
  assign alpha_arctangen_expected_table_data[51] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[52] = 8'b10011111;
  assign alpha_arctangen_expected_table_data[53] = 8'b10100100;
  assign alpha_arctangen_expected_table_data[54] = 8'b10101000;
  assign alpha_arctangen_expected_table_data[55] = 8'b10101100;
  assign alpha_arctangen_expected_table_data[56] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[57] = 8'b10110100;
  assign alpha_arctangen_expected_table_data[58] = 8'b10110010;
  assign alpha_arctangen_expected_table_data[59] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[60] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[61] = 8'b10110011;
  assign alpha_arctangen_expected_table_data[62] = 8'b10111011;
  assign alpha_arctangen_expected_table_data[63] = 8'b11000101;
  assign alpha_arctangen_expected_table_data[64] = 8'b11010110;
  assign alpha_arctangen_expected_table_data[65] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[66] = 8'b11101000;
  assign alpha_arctangen_expected_table_data[67] = 8'b11101100;
  assign alpha_arctangen_expected_table_data[68] = 8'b11101011;
  assign alpha_arctangen_expected_table_data[69] = 8'b11101001;
  assign alpha_arctangen_expected_table_data[70] = 8'b11101000;
  assign alpha_arctangen_expected_table_data[71] = 8'b11101011;
  assign alpha_arctangen_expected_table_data[72] = 8'b11110000;
  assign alpha_arctangen_expected_table_data[73] = 8'b11110100;
  assign alpha_arctangen_expected_table_data[74] = 8'b11111000;
  assign alpha_arctangen_expected_table_data[75] = 8'b11111100;
  assign alpha_arctangen_expected_table_data[76] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[77] = 8'b00000100;
  assign alpha_arctangen_expected_table_data[78] = 8'b00001000;
  assign alpha_arctangen_expected_table_data[79] = 8'b00001100;
  assign alpha_arctangen_expected_table_data[80] = 8'b00010000;
  assign alpha_arctangen_expected_table_data[81] = 8'b00010101;
  assign alpha_arctangen_expected_table_data[82] = 8'b00011000;
  assign alpha_arctangen_expected_table_data[83] = 8'b00010111;
  assign alpha_arctangen_expected_table_data[84] = 8'b00010101;
  assign alpha_arctangen_expected_table_data[85] = 8'b00010100;
  assign alpha_arctangen_expected_table_data[86] = 8'b00011000;
  assign alpha_arctangen_expected_table_data[87] = 8'b00100000;
  assign alpha_arctangen_expected_table_data[88] = 8'b00101010;
  assign alpha_arctangen_expected_table_data[89] = 8'b00111011;
  assign alpha_arctangen_expected_table_data[90] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[91] = 8'b01001101;
  assign alpha_arctangen_expected_table_data[92] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[93] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[94] = 8'b01001110;
  assign alpha_arctangen_expected_table_data[95] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[96] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[97] = 8'b01010100;
  assign alpha_arctangen_expected_table_data[98] = 8'b01011000;
  assign alpha_arctangen_expected_table_data[99] = 8'b01011100;
  assign alpha_arctangen_expected_table_data[100] = 8'b01100001;
  assign alpha_arctangen_expected_table_data[101] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[102] = 8'b10011111;
  assign alpha_arctangen_expected_table_data[103] = 8'b10100100;
  assign alpha_arctangen_expected_table_data[104] = 8'b10101000;
  assign alpha_arctangen_expected_table_data[105] = 8'b10101100;
  assign alpha_arctangen_expected_table_data[106] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[107] = 8'b10110100;
  assign alpha_arctangen_expected_table_data[108] = 8'b10110010;
  assign alpha_arctangen_expected_table_data[109] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[110] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[111] = 8'b10110011;
  assign alpha_arctangen_expected_table_data[112] = 8'b10111011;
  assign alpha_arctangen_expected_table_data[113] = 8'b11000101;
  assign alpha_arctangen_expected_table_data[114] = 8'b11010110;
  assign alpha_arctangen_expected_table_data[115] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[116] = 8'b11101000;
  assign alpha_arctangen_expected_table_data[117] = 8'b11101100;
  assign alpha_arctangen_expected_table_data[118] = 8'b11101011;
  assign alpha_arctangen_expected_table_data[119] = 8'b11101001;
  assign alpha_arctangen_expected_table_data[120] = 8'b11101000;
  assign alpha_arctangen_expected_table_data[121] = 8'b11101011;
  assign alpha_arctangen_expected_table_data[122] = 8'b11110000;
  assign alpha_arctangen_expected_table_data[123] = 8'b11110100;
  assign alpha_arctangen_expected_table_data[124] = 8'b11111000;
  assign alpha_arctangen_expected_table_data[125] = 8'b11111100;
  assign alpha_arctangen_expected_table_data[126] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[127] = 8'b00000100;
  assign alpha_arctangen_expected_table_data[128] = 8'b00001000;
  assign alpha_arctangen_expected_table_data[129] = 8'b00001100;
  assign alpha_arctangen_expected_table_data[130] = 8'b00010000;
  assign alpha_arctangen_expected_table_data[131] = 8'b00010101;
  assign alpha_arctangen_expected_table_data[132] = 8'b00011000;
  assign alpha_arctangen_expected_table_data[133] = 8'b00010111;
  assign alpha_arctangen_expected_table_data[134] = 8'b00010101;
  assign alpha_arctangen_expected_table_data[135] = 8'b00010100;
  assign alpha_arctangen_expected_table_data[136] = 8'b00011000;
  assign alpha_arctangen_expected_table_data[137] = 8'b00100000;
  assign alpha_arctangen_expected_table_data[138] = 8'b00101010;
  assign alpha_arctangen_expected_table_data[139] = 8'b00111011;
  assign alpha_arctangen_expected_table_data[140] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[141] = 8'b01001101;
  assign alpha_arctangen_expected_table_data[142] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[143] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[144] = 8'b01001110;
  assign alpha_arctangen_expected_table_data[145] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[146] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[147] = 8'b01010100;
  assign alpha_arctangen_expected_table_data[148] = 8'b01011000;
  assign alpha_arctangen_expected_table_data[149] = 8'b01011100;
  assign alpha_arctangen_expected_table_data[150] = 8'b01100001;
  assign alpha_arctangen_expected_table_data[151] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[152] = 8'b10011111;
  assign alpha_arctangen_expected_table_data[153] = 8'b10100100;
  assign alpha_arctangen_expected_table_data[154] = 8'b10101000;
  assign alpha_arctangen_expected_table_data[155] = 8'b10101100;
  assign alpha_arctangen_expected_table_data[156] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[157] = 8'b10110100;
  assign alpha_arctangen_expected_table_data[158] = 8'b10110010;
  assign alpha_arctangen_expected_table_data[159] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[160] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[161] = 8'b10110011;
  assign alpha_arctangen_expected_table_data[162] = 8'b10111011;
  assign alpha_arctangen_expected_table_data[163] = 8'b11000101;
  assign alpha_arctangen_expected_table_data[164] = 8'b11010110;
  assign alpha_arctangen_expected_table_data[165] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[166] = 8'b11101000;
  assign alpha_arctangen_expected_table_data[167] = 8'b11101100;
  assign alpha_arctangen_expected_table_data[168] = 8'b11101011;
  assign alpha_arctangen_expected_table_data[169] = 8'b11101001;
  assign alpha_arctangen_expected_table_data[170] = 8'b11101000;
  assign alpha_arctangen_expected_table_data[171] = 8'b11101011;
  assign alpha_arctangen_expected_table_data[172] = 8'b11110000;
  assign alpha_arctangen_expected_table_data[173] = 8'b11110100;
  assign alpha_arctangen_expected_table_data[174] = 8'b11111000;
  assign alpha_arctangen_expected_table_data[175] = 8'b11111100;
  assign alpha_arctangen_expected_table_data[176] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[177] = 8'b00000100;
  assign alpha_arctangen_expected_table_data[178] = 8'b00001000;
  assign alpha_arctangen_expected_table_data[179] = 8'b00001100;
  assign alpha_arctangen_expected_table_data[180] = 8'b00010000;
  assign alpha_arctangen_expected_table_data[181] = 8'b00010101;
  assign alpha_arctangen_expected_table_data[182] = 8'b00011000;
  assign alpha_arctangen_expected_table_data[183] = 8'b00010111;
  assign alpha_arctangen_expected_table_data[184] = 8'b00010101;
  assign alpha_arctangen_expected_table_data[185] = 8'b00010100;
  assign alpha_arctangen_expected_table_data[186] = 8'b00011000;
  assign alpha_arctangen_expected_table_data[187] = 8'b00100000;
  assign alpha_arctangen_expected_table_data[188] = 8'b00101010;
  assign alpha_arctangen_expected_table_data[189] = 8'b00111011;
  assign alpha_arctangen_expected_table_data[190] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[191] = 8'b01001101;
  assign alpha_arctangen_expected_table_data[192] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[193] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[194] = 8'b01001110;
  assign alpha_arctangen_expected_table_data[195] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[196] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[197] = 8'b01010100;
  assign alpha_arctangen_expected_table_data[198] = 8'b01011000;
  assign alpha_arctangen_expected_table_data[199] = 8'b01011100;
  assign alpha_arctangen_expected_table_data[200] = 8'b01100001;
  assign alpha_arctangen_expected_table_data[201] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[202] = 8'b10011111;
  assign alpha_arctangen_expected_table_data[203] = 8'b10100100;
  assign alpha_arctangen_expected_table_data[204] = 8'b10101000;
  assign alpha_arctangen_expected_table_data[205] = 8'b10101100;
  assign alpha_arctangen_expected_table_data[206] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[207] = 8'b10110100;
  assign alpha_arctangen_expected_table_data[208] = 8'b10110010;
  assign alpha_arctangen_expected_table_data[209] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[210] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[211] = 8'b10110011;
  assign alpha_arctangen_expected_table_data[212] = 8'b10111011;
  assign alpha_arctangen_expected_table_data[213] = 8'b11000101;
  assign alpha_arctangen_expected_table_data[214] = 8'b11010110;
  assign alpha_arctangen_expected_table_data[215] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[216] = 8'b11101000;
  assign alpha_arctangen_expected_table_data[217] = 8'b11101100;
  assign alpha_arctangen_expected_table_data[218] = 8'b11101011;
  assign alpha_arctangen_expected_table_data[219] = 8'b11101001;
  assign alpha_arctangen_expected_table_data[220] = 8'b11101000;
  assign alpha_arctangen_expected_table_data[221] = 8'b11101011;
  assign alpha_arctangen_expected_table_data[222] = 8'b11110000;
  assign alpha_arctangen_expected_table_data[223] = 8'b11110100;
  assign alpha_arctangen_expected_table_data[224] = 8'b11111000;
  assign alpha_arctangen_expected_table_data[225] = 8'b11111100;
  assign alpha_arctangen_expected_table_data[226] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[227] = 8'b00000100;
  assign alpha_arctangen_expected_table_data[228] = 8'b00001000;
  assign alpha_arctangen_expected_table_data[229] = 8'b00001100;
  assign alpha_arctangen_expected_table_data[230] = 8'b00010000;
  assign alpha_arctangen_expected_table_data[231] = 8'b00010101;
  assign alpha_arctangen_expected_table_data[232] = 8'b00011000;
  assign alpha_arctangen_expected_table_data[233] = 8'b00010111;
  assign alpha_arctangen_expected_table_data[234] = 8'b00010101;
  assign alpha_arctangen_expected_table_data[235] = 8'b00010100;
  assign alpha_arctangen_expected_table_data[236] = 8'b00011000;
  assign alpha_arctangen_expected_table_data[237] = 8'b00100000;
  assign alpha_arctangen_expected_table_data[238] = 8'b00101010;
  assign alpha_arctangen_expected_table_data[239] = 8'b00111011;
  assign alpha_arctangen_expected_table_data[240] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[241] = 8'b01001101;
  assign alpha_arctangen_expected_table_data[242] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[243] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[244] = 8'b01001110;
  assign alpha_arctangen_expected_table_data[245] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[246] = 8'b01010000;
  assign alpha_arctangen_expected_table_data[247] = 8'b01010100;
  assign alpha_arctangen_expected_table_data[248] = 8'b01011000;
  assign alpha_arctangen_expected_table_data[249] = 8'b01011100;
  assign alpha_arctangen_expected_table_data[250] = 8'b01100001;
  assign alpha_arctangen_expected_table_data[251] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[252] = 8'b10011111;
  assign alpha_arctangen_expected_table_data[253] = 8'b10100100;
  assign alpha_arctangen_expected_table_data[254] = 8'b10101000;
  assign alpha_arctangen_expected_table_data[255] = 8'b10101100;
  assign alpha_arctangen_expected_table_data[256] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[257] = 8'b10110100;
  assign alpha_arctangen_expected_table_data[258] = 8'b10110010;
  assign alpha_arctangen_expected_table_data[259] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[260] = 8'b10110000;
  assign alpha_arctangen_expected_table_data[261] = 8'b10110011;
  assign alpha_arctangen_expected_table_data[262] = 8'b10111011;
  assign alpha_arctangen_expected_table_data[263] = 8'b11000101;
  assign alpha_arctangen_expected_table_data[264] = 8'b11010110;
  assign alpha_arctangen_expected_table_data[265] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[266] = 8'b11101000;
  assign alpha_arctangen_expected_table_data[267] = 8'b11101100;
  assign alpha_arctangen_expected_table_data[268] = 8'b11101011;
  assign alpha_arctangen_expected_table_data[269] = 8'b11101001;
  assign alpha_arctangen_expected_table_data[270] = 8'b11101000;
  assign alpha_arctangen_expected_table_data[271] = 8'b11101011;
  assign alpha_arctangen_expected_table_data[272] = 8'b11110000;
  assign alpha_arctangen_expected_table_data[273] = 8'b11110100;
  assign alpha_arctangen_expected_table_data[274] = 8'b11111000;
  assign alpha_arctangen_expected_table_data[275] = 8'b11111100;
  assign alpha_arctangen_expected_table_data[276] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[277] = 8'b10100000;
  assign alpha_arctangen_expected_table_data[278] = 8'b10100011;
  assign alpha_arctangen_expected_table_data[279] = 8'b10100101;
  assign alpha_arctangen_expected_table_data[280] = 8'b10101010;
  assign alpha_arctangen_expected_table_data[281] = 8'b10101011;
  assign alpha_arctangen_expected_table_data[282] = 8'b10101101;
  assign alpha_arctangen_expected_table_data[283] = 8'b10111100;
  assign alpha_arctangen_expected_table_data[284] = 8'b10111011;
  assign alpha_arctangen_expected_table_data[285] = 8'b10111110;
  assign alpha_arctangen_expected_table_data[286] = 8'b11000000;
  assign alpha_arctangen_expected_table_data[287] = 8'b11000111;
  assign alpha_arctangen_expected_table_data[288] = 8'b11001010;
  assign alpha_arctangen_expected_table_data[289] = 8'b11010001;
  assign alpha_arctangen_expected_table_data[290] = 8'b11010101;
  assign alpha_arctangen_expected_table_data[291] = 8'b11011011;
  assign alpha_arctangen_expected_table_data[292] = 8'b11011101;
  assign alpha_arctangen_expected_table_data[293] = 8'b11100001;
  assign alpha_arctangen_expected_table_data[294] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[295] = 8'b11101110;
  assign alpha_arctangen_expected_table_data[296] = 8'b11110000;
  assign alpha_arctangen_expected_table_data[297] = 8'b11110010;
  assign alpha_arctangen_expected_table_data[298] = 8'b11110110;
  assign alpha_arctangen_expected_table_data[299] = 8'b11111000;
  assign alpha_arctangen_expected_table_data[300] = 8'b11111100;
  assign alpha_arctangen_expected_table_data[301] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[302] = 8'b00000100;
  assign alpha_arctangen_expected_table_data[303] = 8'b00001000;
  assign alpha_arctangen_expected_table_data[304] = 8'b00001010;
  assign alpha_arctangen_expected_table_data[305] = 8'b00001110;
  assign alpha_arctangen_expected_table_data[306] = 8'b00010000;
  assign alpha_arctangen_expected_table_data[307] = 8'b00010010;
  assign alpha_arctangen_expected_table_data[308] = 8'b00100000;
  assign alpha_arctangen_expected_table_data[309] = 8'b00011111;
  assign alpha_arctangen_expected_table_data[310] = 8'b00100011;
  assign alpha_arctangen_expected_table_data[311] = 8'b00100101;
  assign alpha_arctangen_expected_table_data[312] = 8'b00101011;
  assign alpha_arctangen_expected_table_data[313] = 8'b00101111;
  assign alpha_arctangen_expected_table_data[314] = 8'b00110110;
  assign alpha_arctangen_expected_table_data[315] = 8'b00111001;
  assign alpha_arctangen_expected_table_data[316] = 8'b01000000;
  assign alpha_arctangen_expected_table_data[317] = 8'b01000010;
  assign alpha_arctangen_expected_table_data[318] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[319] = 8'b01000100;
  assign alpha_arctangen_expected_table_data[320] = 8'b01010011;
  assign alpha_arctangen_expected_table_data[321] = 8'b01010101;
  assign alpha_arctangen_expected_table_data[322] = 8'b01010110;
  assign alpha_arctangen_expected_table_data[323] = 8'b01011011;
  assign alpha_arctangen_expected_table_data[324] = 8'b01011101;
  assign alpha_arctangen_expected_table_data[325] = 8'b01100000;
  assign alpha_arctangen_expected_table_data[326] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[327] = 8'b10100000;
  assign alpha_arctangen_expected_table_data[328] = 8'b10100011;
  assign alpha_arctangen_expected_table_data[329] = 8'b10100101;
  assign alpha_arctangen_expected_table_data[330] = 8'b10101010;
  assign alpha_arctangen_expected_table_data[331] = 8'b10101011;
  assign alpha_arctangen_expected_table_data[332] = 8'b10101101;
  assign alpha_arctangen_expected_table_data[333] = 8'b10111100;
  assign alpha_arctangen_expected_table_data[334] = 8'b10111011;
  assign alpha_arctangen_expected_table_data[335] = 8'b10111110;
  assign alpha_arctangen_expected_table_data[336] = 8'b11000000;
  assign alpha_arctangen_expected_table_data[337] = 8'b11000111;
  assign alpha_arctangen_expected_table_data[338] = 8'b11001010;
  assign alpha_arctangen_expected_table_data[339] = 8'b11010001;
  assign alpha_arctangen_expected_table_data[340] = 8'b11010101;
  assign alpha_arctangen_expected_table_data[341] = 8'b11011011;
  assign alpha_arctangen_expected_table_data[342] = 8'b11011101;
  assign alpha_arctangen_expected_table_data[343] = 8'b11100001;
  assign alpha_arctangen_expected_table_data[344] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[345] = 8'b11101110;
  assign alpha_arctangen_expected_table_data[346] = 8'b11110000;
  assign alpha_arctangen_expected_table_data[347] = 8'b11110010;
  assign alpha_arctangen_expected_table_data[348] = 8'b11110110;
  assign alpha_arctangen_expected_table_data[349] = 8'b11111000;
  assign alpha_arctangen_expected_table_data[350] = 8'b11111100;
  assign alpha_arctangen_expected_table_data[351] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[352] = 8'b00000100;
  assign alpha_arctangen_expected_table_data[353] = 8'b00001000;
  assign alpha_arctangen_expected_table_data[354] = 8'b00001010;
  assign alpha_arctangen_expected_table_data[355] = 8'b00001110;
  assign alpha_arctangen_expected_table_data[356] = 8'b00010000;
  assign alpha_arctangen_expected_table_data[357] = 8'b00010010;
  assign alpha_arctangen_expected_table_data[358] = 8'b00100000;
  assign alpha_arctangen_expected_table_data[359] = 8'b00011111;
  assign alpha_arctangen_expected_table_data[360] = 8'b00100011;
  assign alpha_arctangen_expected_table_data[361] = 8'b00100101;
  assign alpha_arctangen_expected_table_data[362] = 8'b00101011;
  assign alpha_arctangen_expected_table_data[363] = 8'b00101111;
  assign alpha_arctangen_expected_table_data[364] = 8'b00110110;
  assign alpha_arctangen_expected_table_data[365] = 8'b00111001;
  assign alpha_arctangen_expected_table_data[366] = 8'b01000000;
  assign alpha_arctangen_expected_table_data[367] = 8'b01000010;
  assign alpha_arctangen_expected_table_data[368] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[369] = 8'b01000100;
  assign alpha_arctangen_expected_table_data[370] = 8'b01010011;
  assign alpha_arctangen_expected_table_data[371] = 8'b01010101;
  assign alpha_arctangen_expected_table_data[372] = 8'b01010110;
  assign alpha_arctangen_expected_table_data[373] = 8'b01011011;
  assign alpha_arctangen_expected_table_data[374] = 8'b01011101;
  assign alpha_arctangen_expected_table_data[375] = 8'b01100000;
  assign alpha_arctangen_expected_table_data[376] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[377] = 8'b10100000;
  assign alpha_arctangen_expected_table_data[378] = 8'b10100011;
  assign alpha_arctangen_expected_table_data[379] = 8'b10100101;
  assign alpha_arctangen_expected_table_data[380] = 8'b10101010;
  assign alpha_arctangen_expected_table_data[381] = 8'b10101011;
  assign alpha_arctangen_expected_table_data[382] = 8'b10101101;
  assign alpha_arctangen_expected_table_data[383] = 8'b10111100;
  assign alpha_arctangen_expected_table_data[384] = 8'b10111011;
  assign alpha_arctangen_expected_table_data[385] = 8'b10111110;
  assign alpha_arctangen_expected_table_data[386] = 8'b11000000;
  assign alpha_arctangen_expected_table_data[387] = 8'b11000111;
  assign alpha_arctangen_expected_table_data[388] = 8'b11001010;
  assign alpha_arctangen_expected_table_data[389] = 8'b11010001;
  assign alpha_arctangen_expected_table_data[390] = 8'b11010101;
  assign alpha_arctangen_expected_table_data[391] = 8'b11011011;
  assign alpha_arctangen_expected_table_data[392] = 8'b11011101;
  assign alpha_arctangen_expected_table_data[393] = 8'b11100001;
  assign alpha_arctangen_expected_table_data[394] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[395] = 8'b11101110;
  assign alpha_arctangen_expected_table_data[396] = 8'b11110000;
  assign alpha_arctangen_expected_table_data[397] = 8'b11110010;
  assign alpha_arctangen_expected_table_data[398] = 8'b11110110;
  assign alpha_arctangen_expected_table_data[399] = 8'b11111000;
  assign alpha_arctangen_expected_table_data[400] = 8'b11111100;
  assign alpha_arctangen_expected_table_data[401] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[402] = 8'b00000100;
  assign alpha_arctangen_expected_table_data[403] = 8'b00001000;
  assign alpha_arctangen_expected_table_data[404] = 8'b00001010;
  assign alpha_arctangen_expected_table_data[405] = 8'b00001110;
  assign alpha_arctangen_expected_table_data[406] = 8'b00010000;
  assign alpha_arctangen_expected_table_data[407] = 8'b00010010;
  assign alpha_arctangen_expected_table_data[408] = 8'b00100000;
  assign alpha_arctangen_expected_table_data[409] = 8'b00011111;
  assign alpha_arctangen_expected_table_data[410] = 8'b00100011;
  assign alpha_arctangen_expected_table_data[411] = 8'b00100101;
  assign alpha_arctangen_expected_table_data[412] = 8'b00101011;
  assign alpha_arctangen_expected_table_data[413] = 8'b00101111;
  assign alpha_arctangen_expected_table_data[414] = 8'b00110110;
  assign alpha_arctangen_expected_table_data[415] = 8'b00111001;
  assign alpha_arctangen_expected_table_data[416] = 8'b01000000;
  assign alpha_arctangen_expected_table_data[417] = 8'b01000010;
  assign alpha_arctangen_expected_table_data[418] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[419] = 8'b01000100;
  assign alpha_arctangen_expected_table_data[420] = 8'b01010011;
  assign alpha_arctangen_expected_table_data[421] = 8'b01010101;
  assign alpha_arctangen_expected_table_data[422] = 8'b01010110;
  assign alpha_arctangen_expected_table_data[423] = 8'b01011011;
  assign alpha_arctangen_expected_table_data[424] = 8'b01011101;
  assign alpha_arctangen_expected_table_data[425] = 8'b01100000;
  assign alpha_arctangen_expected_table_data[426] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[427] = 8'b10100000;
  assign alpha_arctangen_expected_table_data[428] = 8'b10100011;
  assign alpha_arctangen_expected_table_data[429] = 8'b10100101;
  assign alpha_arctangen_expected_table_data[430] = 8'b10101010;
  assign alpha_arctangen_expected_table_data[431] = 8'b10101011;
  assign alpha_arctangen_expected_table_data[432] = 8'b10101101;
  assign alpha_arctangen_expected_table_data[433] = 8'b10111100;
  assign alpha_arctangen_expected_table_data[434] = 8'b10111011;
  assign alpha_arctangen_expected_table_data[435] = 8'b10111110;
  assign alpha_arctangen_expected_table_data[436] = 8'b11000000;
  assign alpha_arctangen_expected_table_data[437] = 8'b11000111;
  assign alpha_arctangen_expected_table_data[438] = 8'b11001010;
  assign alpha_arctangen_expected_table_data[439] = 8'b11010001;
  assign alpha_arctangen_expected_table_data[440] = 8'b11010101;
  assign alpha_arctangen_expected_table_data[441] = 8'b11011011;
  assign alpha_arctangen_expected_table_data[442] = 8'b11011101;
  assign alpha_arctangen_expected_table_data[443] = 8'b11100001;
  assign alpha_arctangen_expected_table_data[444] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[445] = 8'b11101110;
  assign alpha_arctangen_expected_table_data[446] = 8'b11110000;
  assign alpha_arctangen_expected_table_data[447] = 8'b11110010;
  assign alpha_arctangen_expected_table_data[448] = 8'b11110110;
  assign alpha_arctangen_expected_table_data[449] = 8'b11111000;
  assign alpha_arctangen_expected_table_data[450] = 8'b11111100;
  assign alpha_arctangen_expected_table_data[451] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[452] = 8'b00000100;
  assign alpha_arctangen_expected_table_data[453] = 8'b00001000;
  assign alpha_arctangen_expected_table_data[454] = 8'b00001010;
  assign alpha_arctangen_expected_table_data[455] = 8'b00001110;
  assign alpha_arctangen_expected_table_data[456] = 8'b00010000;
  assign alpha_arctangen_expected_table_data[457] = 8'b00010010;
  assign alpha_arctangen_expected_table_data[458] = 8'b00100000;
  assign alpha_arctangen_expected_table_data[459] = 8'b00011111;
  assign alpha_arctangen_expected_table_data[460] = 8'b00100011;
  assign alpha_arctangen_expected_table_data[461] = 8'b00100101;
  assign alpha_arctangen_expected_table_data[462] = 8'b00101011;
  assign alpha_arctangen_expected_table_data[463] = 8'b00101111;
  assign alpha_arctangen_expected_table_data[464] = 8'b00110110;
  assign alpha_arctangen_expected_table_data[465] = 8'b00111001;
  assign alpha_arctangen_expected_table_data[466] = 8'b01000000;
  assign alpha_arctangen_expected_table_data[467] = 8'b01000010;
  assign alpha_arctangen_expected_table_data[468] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[469] = 8'b01000100;
  assign alpha_arctangen_expected_table_data[470] = 8'b01010011;
  assign alpha_arctangen_expected_table_data[471] = 8'b01010101;
  assign alpha_arctangen_expected_table_data[472] = 8'b01010110;
  assign alpha_arctangen_expected_table_data[473] = 8'b01011011;
  assign alpha_arctangen_expected_table_data[474] = 8'b01011101;
  assign alpha_arctangen_expected_table_data[475] = 8'b01100000;
  assign alpha_arctangen_expected_table_data[476] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[477] = 8'b10100000;
  assign alpha_arctangen_expected_table_data[478] = 8'b10100011;
  assign alpha_arctangen_expected_table_data[479] = 8'b10100101;
  assign alpha_arctangen_expected_table_data[480] = 8'b10101010;
  assign alpha_arctangen_expected_table_data[481] = 8'b10101011;
  assign alpha_arctangen_expected_table_data[482] = 8'b10101101;
  assign alpha_arctangen_expected_table_data[483] = 8'b10111100;
  assign alpha_arctangen_expected_table_data[484] = 8'b10111011;
  assign alpha_arctangen_expected_table_data[485] = 8'b10111110;
  assign alpha_arctangen_expected_table_data[486] = 8'b11000000;
  assign alpha_arctangen_expected_table_data[487] = 8'b11000111;
  assign alpha_arctangen_expected_table_data[488] = 8'b11001010;
  assign alpha_arctangen_expected_table_data[489] = 8'b11010001;
  assign alpha_arctangen_expected_table_data[490] = 8'b11010101;
  assign alpha_arctangen_expected_table_data[491] = 8'b11011011;
  assign alpha_arctangen_expected_table_data[492] = 8'b11011101;
  assign alpha_arctangen_expected_table_data[493] = 8'b11100001;
  assign alpha_arctangen_expected_table_data[494] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[495] = 8'b11101110;
  assign alpha_arctangen_expected_table_data[496] = 8'b11110000;
  assign alpha_arctangen_expected_table_data[497] = 8'b11110010;
  assign alpha_arctangen_expected_table_data[498] = 8'b11110110;
  assign alpha_arctangen_expected_table_data[499] = 8'b11111000;
  assign alpha_arctangen_expected_table_data[500] = 8'b11111100;
  assign alpha_arctangen_expected_table_data[501] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[502] = 8'b00000100;
  assign alpha_arctangen_expected_table_data[503] = 8'b00001000;
  assign alpha_arctangen_expected_table_data[504] = 8'b00001010;
  assign alpha_arctangen_expected_table_data[505] = 8'b00001110;
  assign alpha_arctangen_expected_table_data[506] = 8'b00010000;
  assign alpha_arctangen_expected_table_data[507] = 8'b00010010;
  assign alpha_arctangen_expected_table_data[508] = 8'b00100000;
  assign alpha_arctangen_expected_table_data[509] = 8'b00011111;
  assign alpha_arctangen_expected_table_data[510] = 8'b00100011;
  assign alpha_arctangen_expected_table_data[511] = 8'b00100101;
  assign alpha_arctangen_expected_table_data[512] = 8'b00101011;
  assign alpha_arctangen_expected_table_data[513] = 8'b00101111;
  assign alpha_arctangen_expected_table_data[514] = 8'b00110110;
  assign alpha_arctangen_expected_table_data[515] = 8'b00111001;
  assign alpha_arctangen_expected_table_data[516] = 8'b01000000;
  assign alpha_arctangen_expected_table_data[517] = 8'b01000010;
  assign alpha_arctangen_expected_table_data[518] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[519] = 8'b01000100;
  assign alpha_arctangen_expected_table_data[520] = 8'b01010011;
  assign alpha_arctangen_expected_table_data[521] = 8'b01010101;
  assign alpha_arctangen_expected_table_data[522] = 8'b01010110;
  assign alpha_arctangen_expected_table_data[523] = 8'b01011011;
  assign alpha_arctangen_expected_table_data[524] = 8'b01011101;
  assign alpha_arctangen_expected_table_data[525] = 8'b01100000;
  assign alpha_arctangen_expected_table_data[526] = 8'b11100111;
  assign alpha_arctangen_expected_table_data[527] = 8'b11100111;
  assign alpha_arctangen_expected_table_data[528] = 8'b11101001;
  assign alpha_arctangen_expected_table_data[529] = 8'b11101100;
  assign alpha_arctangen_expected_table_data[530] = 8'b11101111;
  assign alpha_arctangen_expected_table_data[531] = 8'b11110010;
  assign alpha_arctangen_expected_table_data[532] = 8'b11110110;
  assign alpha_arctangen_expected_table_data[533] = 8'b11111010;
  assign alpha_arctangen_expected_table_data[534] = 8'b11111111;
  assign alpha_arctangen_expected_table_data[535] = 8'b00000010;
  assign alpha_arctangen_expected_table_data[536] = 8'b00000111;
  assign alpha_arctangen_expected_table_data[537] = 8'b00001011;
  assign alpha_arctangen_expected_table_data[538] = 8'b00001111;
  assign alpha_arctangen_expected_table_data[539] = 8'b00010010;
  assign alpha_arctangen_expected_table_data[540] = 8'b00010110;
  assign alpha_arctangen_expected_table_data[541] = 8'b00011001;
  assign alpha_arctangen_expected_table_data[542] = 8'b00011001;
  assign alpha_arctangen_expected_table_data[543] = 8'b00011010;
  assign alpha_arctangen_expected_table_data[544] = 8'b00011101;
  assign alpha_arctangen_expected_table_data[545] = 8'b00100011;
  assign alpha_arctangen_expected_table_data[546] = 8'b00101010;
  assign alpha_arctangen_expected_table_data[547] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[548] = 8'b00111111;
  assign alpha_arctangen_expected_table_data[549] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[550] = 8'b01001010;
  assign alpha_arctangen_expected_table_data[551] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[552] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[553] = 8'b01001101;
  assign alpha_arctangen_expected_table_data[554] = 8'b01010001;
  assign alpha_arctangen_expected_table_data[555] = 8'b01010100;
  assign alpha_arctangen_expected_table_data[556] = 8'b01010111;
  assign alpha_arctangen_expected_table_data[557] = 8'b01011010;
  assign alpha_arctangen_expected_table_data[558] = 8'b01011111;
  assign alpha_arctangen_expected_table_data[559] = 8'b01100011;
  assign alpha_arctangen_expected_table_data[560] = 8'b10011110;
  assign alpha_arctangen_expected_table_data[561] = 8'b10100010;
  assign alpha_arctangen_expected_table_data[562] = 8'b10100111;
  assign alpha_arctangen_expected_table_data[563] = 8'b10101010;
  assign alpha_arctangen_expected_table_data[564] = 8'b10101110;
  assign alpha_arctangen_expected_table_data[565] = 8'b10110001;
  assign alpha_arctangen_expected_table_data[566] = 8'b10110101;
  assign alpha_arctangen_expected_table_data[567] = 8'b10110100;
  assign alpha_arctangen_expected_table_data[568] = 8'b10110101;
  assign alpha_arctangen_expected_table_data[569] = 8'b10111000;
  assign alpha_arctangen_expected_table_data[570] = 8'b10111110;
  assign alpha_arctangen_expected_table_data[571] = 8'b11000101;
  assign alpha_arctangen_expected_table_data[572] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[573] = 8'b11011010;
  assign alpha_arctangen_expected_table_data[574] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[575] = 8'b11100101;
  assign alpha_arctangen_expected_table_data[576] = 8'b11100111;
  assign alpha_arctangen_expected_table_data[577] = 8'b11100111;
  assign alpha_arctangen_expected_table_data[578] = 8'b11101001;
  assign alpha_arctangen_expected_table_data[579] = 8'b11101100;
  assign alpha_arctangen_expected_table_data[580] = 8'b11101111;
  assign alpha_arctangen_expected_table_data[581] = 8'b11110010;
  assign alpha_arctangen_expected_table_data[582] = 8'b11110110;
  assign alpha_arctangen_expected_table_data[583] = 8'b11111010;
  assign alpha_arctangen_expected_table_data[584] = 8'b11111111;
  assign alpha_arctangen_expected_table_data[585] = 8'b00000010;
  assign alpha_arctangen_expected_table_data[586] = 8'b00000111;
  assign alpha_arctangen_expected_table_data[587] = 8'b00001011;
  assign alpha_arctangen_expected_table_data[588] = 8'b00001111;
  assign alpha_arctangen_expected_table_data[589] = 8'b00010010;
  assign alpha_arctangen_expected_table_data[590] = 8'b00010110;
  assign alpha_arctangen_expected_table_data[591] = 8'b00011001;
  assign alpha_arctangen_expected_table_data[592] = 8'b00011001;
  assign alpha_arctangen_expected_table_data[593] = 8'b00011010;
  assign alpha_arctangen_expected_table_data[594] = 8'b00011101;
  assign alpha_arctangen_expected_table_data[595] = 8'b00100011;
  assign alpha_arctangen_expected_table_data[596] = 8'b00101010;
  assign alpha_arctangen_expected_table_data[597] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[598] = 8'b00111111;
  assign alpha_arctangen_expected_table_data[599] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[600] = 8'b01001010;
  assign alpha_arctangen_expected_table_data[601] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[602] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[603] = 8'b01001101;
  assign alpha_arctangen_expected_table_data[604] = 8'b01010001;
  assign alpha_arctangen_expected_table_data[605] = 8'b01010100;
  assign alpha_arctangen_expected_table_data[606] = 8'b01010111;
  assign alpha_arctangen_expected_table_data[607] = 8'b01011010;
  assign alpha_arctangen_expected_table_data[608] = 8'b01011111;
  assign alpha_arctangen_expected_table_data[609] = 8'b01100011;
  assign alpha_arctangen_expected_table_data[610] = 8'b10011110;
  assign alpha_arctangen_expected_table_data[611] = 8'b10100010;
  assign alpha_arctangen_expected_table_data[612] = 8'b10100111;
  assign alpha_arctangen_expected_table_data[613] = 8'b10101010;
  assign alpha_arctangen_expected_table_data[614] = 8'b10101110;
  assign alpha_arctangen_expected_table_data[615] = 8'b10110001;
  assign alpha_arctangen_expected_table_data[616] = 8'b10110101;
  assign alpha_arctangen_expected_table_data[617] = 8'b10110100;
  assign alpha_arctangen_expected_table_data[618] = 8'b10110101;
  assign alpha_arctangen_expected_table_data[619] = 8'b10111000;
  assign alpha_arctangen_expected_table_data[620] = 8'b10111110;
  assign alpha_arctangen_expected_table_data[621] = 8'b11000101;
  assign alpha_arctangen_expected_table_data[622] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[623] = 8'b11011010;
  assign alpha_arctangen_expected_table_data[624] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[625] = 8'b11100101;
  assign alpha_arctangen_expected_table_data[626] = 8'b11100111;
  assign alpha_arctangen_expected_table_data[627] = 8'b11100111;
  assign alpha_arctangen_expected_table_data[628] = 8'b11101001;
  assign alpha_arctangen_expected_table_data[629] = 8'b11101100;
  assign alpha_arctangen_expected_table_data[630] = 8'b11101111;
  assign alpha_arctangen_expected_table_data[631] = 8'b11110010;
  assign alpha_arctangen_expected_table_data[632] = 8'b11110110;
  assign alpha_arctangen_expected_table_data[633] = 8'b11111010;
  assign alpha_arctangen_expected_table_data[634] = 8'b11111111;
  assign alpha_arctangen_expected_table_data[635] = 8'b00000010;
  assign alpha_arctangen_expected_table_data[636] = 8'b00000111;
  assign alpha_arctangen_expected_table_data[637] = 8'b00001011;
  assign alpha_arctangen_expected_table_data[638] = 8'b00001111;
  assign alpha_arctangen_expected_table_data[639] = 8'b00010010;
  assign alpha_arctangen_expected_table_data[640] = 8'b00010110;
  assign alpha_arctangen_expected_table_data[641] = 8'b00011001;
  assign alpha_arctangen_expected_table_data[642] = 8'b00011001;
  assign alpha_arctangen_expected_table_data[643] = 8'b00011010;
  assign alpha_arctangen_expected_table_data[644] = 8'b00011101;
  assign alpha_arctangen_expected_table_data[645] = 8'b00100011;
  assign alpha_arctangen_expected_table_data[646] = 8'b00101010;
  assign alpha_arctangen_expected_table_data[647] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[648] = 8'b00111111;
  assign alpha_arctangen_expected_table_data[649] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[650] = 8'b01001010;
  assign alpha_arctangen_expected_table_data[651] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[652] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[653] = 8'b01001101;
  assign alpha_arctangen_expected_table_data[654] = 8'b01010001;
  assign alpha_arctangen_expected_table_data[655] = 8'b01010100;
  assign alpha_arctangen_expected_table_data[656] = 8'b01010111;
  assign alpha_arctangen_expected_table_data[657] = 8'b01011010;
  assign alpha_arctangen_expected_table_data[658] = 8'b01011111;
  assign alpha_arctangen_expected_table_data[659] = 8'b01100011;
  assign alpha_arctangen_expected_table_data[660] = 8'b10011110;
  assign alpha_arctangen_expected_table_data[661] = 8'b10100010;
  assign alpha_arctangen_expected_table_data[662] = 8'b10100111;
  assign alpha_arctangen_expected_table_data[663] = 8'b10101010;
  assign alpha_arctangen_expected_table_data[664] = 8'b10101110;
  assign alpha_arctangen_expected_table_data[665] = 8'b10110001;
  assign alpha_arctangen_expected_table_data[666] = 8'b10110101;
  assign alpha_arctangen_expected_table_data[667] = 8'b10110100;
  assign alpha_arctangen_expected_table_data[668] = 8'b10110101;
  assign alpha_arctangen_expected_table_data[669] = 8'b10111000;
  assign alpha_arctangen_expected_table_data[670] = 8'b10111110;
  assign alpha_arctangen_expected_table_data[671] = 8'b11000101;
  assign alpha_arctangen_expected_table_data[672] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[673] = 8'b11011010;
  assign alpha_arctangen_expected_table_data[674] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[675] = 8'b11100101;
  assign alpha_arctangen_expected_table_data[676] = 8'b11100111;
  assign alpha_arctangen_expected_table_data[677] = 8'b11100111;
  assign alpha_arctangen_expected_table_data[678] = 8'b11101001;
  assign alpha_arctangen_expected_table_data[679] = 8'b11101100;
  assign alpha_arctangen_expected_table_data[680] = 8'b11101111;
  assign alpha_arctangen_expected_table_data[681] = 8'b11110010;
  assign alpha_arctangen_expected_table_data[682] = 8'b11110110;
  assign alpha_arctangen_expected_table_data[683] = 8'b11111010;
  assign alpha_arctangen_expected_table_data[684] = 8'b11111111;
  assign alpha_arctangen_expected_table_data[685] = 8'b00000010;
  assign alpha_arctangen_expected_table_data[686] = 8'b00000111;
  assign alpha_arctangen_expected_table_data[687] = 8'b00001011;
  assign alpha_arctangen_expected_table_data[688] = 8'b00001111;
  assign alpha_arctangen_expected_table_data[689] = 8'b00010010;
  assign alpha_arctangen_expected_table_data[690] = 8'b00010110;
  assign alpha_arctangen_expected_table_data[691] = 8'b00011001;
  assign alpha_arctangen_expected_table_data[692] = 8'b00011001;
  assign alpha_arctangen_expected_table_data[693] = 8'b00011010;
  assign alpha_arctangen_expected_table_data[694] = 8'b00011101;
  assign alpha_arctangen_expected_table_data[695] = 8'b00100011;
  assign alpha_arctangen_expected_table_data[696] = 8'b00101010;
  assign alpha_arctangen_expected_table_data[697] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[698] = 8'b00111111;
  assign alpha_arctangen_expected_table_data[699] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[700] = 8'b01001010;
  assign alpha_arctangen_expected_table_data[701] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[702] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[703] = 8'b01001101;
  assign alpha_arctangen_expected_table_data[704] = 8'b01010001;
  assign alpha_arctangen_expected_table_data[705] = 8'b01010100;
  assign alpha_arctangen_expected_table_data[706] = 8'b01010111;
  assign alpha_arctangen_expected_table_data[707] = 8'b01011010;
  assign alpha_arctangen_expected_table_data[708] = 8'b01011111;
  assign alpha_arctangen_expected_table_data[709] = 8'b01100011;
  assign alpha_arctangen_expected_table_data[710] = 8'b10011110;
  assign alpha_arctangen_expected_table_data[711] = 8'b10100010;
  assign alpha_arctangen_expected_table_data[712] = 8'b10100111;
  assign alpha_arctangen_expected_table_data[713] = 8'b10101010;
  assign alpha_arctangen_expected_table_data[714] = 8'b10101110;
  assign alpha_arctangen_expected_table_data[715] = 8'b10110001;
  assign alpha_arctangen_expected_table_data[716] = 8'b10110101;
  assign alpha_arctangen_expected_table_data[717] = 8'b10110100;
  assign alpha_arctangen_expected_table_data[718] = 8'b10110101;
  assign alpha_arctangen_expected_table_data[719] = 8'b10111000;
  assign alpha_arctangen_expected_table_data[720] = 8'b10111110;
  assign alpha_arctangen_expected_table_data[721] = 8'b11000101;
  assign alpha_arctangen_expected_table_data[722] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[723] = 8'b11011010;
  assign alpha_arctangen_expected_table_data[724] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[725] = 8'b11100101;
  assign alpha_arctangen_expected_table_data[726] = 8'b11100111;
  assign alpha_arctangen_expected_table_data[727] = 8'b11100111;
  assign alpha_arctangen_expected_table_data[728] = 8'b11101001;
  assign alpha_arctangen_expected_table_data[729] = 8'b11101100;
  assign alpha_arctangen_expected_table_data[730] = 8'b11101111;
  assign alpha_arctangen_expected_table_data[731] = 8'b11110010;
  assign alpha_arctangen_expected_table_data[732] = 8'b11110110;
  assign alpha_arctangen_expected_table_data[733] = 8'b11111010;
  assign alpha_arctangen_expected_table_data[734] = 8'b11111111;
  assign alpha_arctangen_expected_table_data[735] = 8'b00000010;
  assign alpha_arctangen_expected_table_data[736] = 8'b00000111;
  assign alpha_arctangen_expected_table_data[737] = 8'b00001011;
  assign alpha_arctangen_expected_table_data[738] = 8'b00001111;
  assign alpha_arctangen_expected_table_data[739] = 8'b00010010;
  assign alpha_arctangen_expected_table_data[740] = 8'b00010110;
  assign alpha_arctangen_expected_table_data[741] = 8'b00011001;
  assign alpha_arctangen_expected_table_data[742] = 8'b00011001;
  assign alpha_arctangen_expected_table_data[743] = 8'b00011010;
  assign alpha_arctangen_expected_table_data[744] = 8'b00011101;
  assign alpha_arctangen_expected_table_data[745] = 8'b00100011;
  assign alpha_arctangen_expected_table_data[746] = 8'b00101010;
  assign alpha_arctangen_expected_table_data[747] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[748] = 8'b00111111;
  assign alpha_arctangen_expected_table_data[749] = 8'b01000101;
  assign alpha_arctangen_expected_table_data[750] = 8'b01001010;
  assign alpha_arctangen_expected_table_data[751] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[752] = 8'b01001100;
  assign alpha_arctangen_expected_table_data[753] = 8'b01001101;
  assign alpha_arctangen_expected_table_data[754] = 8'b01010001;
  assign alpha_arctangen_expected_table_data[755] = 8'b01010100;
  assign alpha_arctangen_expected_table_data[756] = 8'b01010111;
  assign alpha_arctangen_expected_table_data[757] = 8'b01011010;
  assign alpha_arctangen_expected_table_data[758] = 8'b01011111;
  assign alpha_arctangen_expected_table_data[759] = 8'b01100011;
  assign alpha_arctangen_expected_table_data[760] = 8'b10011110;
  assign alpha_arctangen_expected_table_data[761] = 8'b10100010;
  assign alpha_arctangen_expected_table_data[762] = 8'b10100111;
  assign alpha_arctangen_expected_table_data[763] = 8'b10101010;
  assign alpha_arctangen_expected_table_data[764] = 8'b10101110;
  assign alpha_arctangen_expected_table_data[765] = 8'b10110001;
  assign alpha_arctangen_expected_table_data[766] = 8'b10110101;
  assign alpha_arctangen_expected_table_data[767] = 8'b10110100;
  assign alpha_arctangen_expected_table_data[768] = 8'b10110101;
  assign alpha_arctangen_expected_table_data[769] = 8'b10111000;
  assign alpha_arctangen_expected_table_data[770] = 8'b10111110;
  assign alpha_arctangen_expected_table_data[771] = 8'b11000101;
  assign alpha_arctangen_expected_table_data[772] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[773] = 8'b11011010;
  assign alpha_arctangen_expected_table_data[774] = 8'b11100000;
  assign alpha_arctangen_expected_table_data[775] = 8'b11100101;
  assign alpha_arctangen_expected_table_data[776] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[777] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[778] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[779] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[780] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[781] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[782] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[783] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[784] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[785] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[786] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[787] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[788] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[789] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[790] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[791] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[792] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[793] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[794] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[795] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[796] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[797] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[798] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[799] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[800] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[801] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[802] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[803] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[804] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[805] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[806] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[807] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[808] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[809] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[810] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[811] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[812] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[813] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[814] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[815] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[816] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[817] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[818] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[819] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[820] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[821] = 8'b11111111;
  assign alpha_arctangen_expected_table_data[822] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[823] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[824] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[825] = 8'b00000001;
  assign alpha_arctangen_expected_table_data[826] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[827] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[828] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[829] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[830] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[831] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[832] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[833] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[834] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[835] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[836] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[837] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[838] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[839] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[840] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[841] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[842] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[843] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[844] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[845] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[846] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[847] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[848] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[849] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[850] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[851] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[852] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[853] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[854] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[855] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[856] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[857] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[858] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[859] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[860] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[861] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[862] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[863] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[864] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[865] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[866] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[867] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[868] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[869] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[870] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[871] = 8'b11111111;
  assign alpha_arctangen_expected_table_data[872] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[873] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[874] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[875] = 8'b00000001;
  assign alpha_arctangen_expected_table_data[876] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[877] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[878] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[879] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[880] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[881] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[882] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[883] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[884] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[885] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[886] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[887] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[888] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[889] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[890] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[891] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[892] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[893] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[894] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[895] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[896] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[897] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[898] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[899] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[900] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[901] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[902] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[903] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[904] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[905] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[906] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[907] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[908] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[909] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[910] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[911] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[912] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[913] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[914] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[915] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[916] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[917] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[918] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[919] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[920] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[921] = 8'b11111111;
  assign alpha_arctangen_expected_table_data[922] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[923] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[924] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[925] = 8'b00000001;
  assign alpha_arctangen_expected_table_data[926] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[927] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[928] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[929] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[930] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[931] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[932] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[933] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[934] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[935] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[936] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[937] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[938] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[939] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[940] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[941] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[942] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[943] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[944] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[945] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[946] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[947] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[948] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[949] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[950] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[951] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[952] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[953] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[954] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[955] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[956] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[957] = 8'b11001101;
  assign alpha_arctangen_expected_table_data[958] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[959] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[960] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[961] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[962] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[963] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[964] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[965] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[966] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[967] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[968] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[969] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[970] = 8'b11001110;
  assign alpha_arctangen_expected_table_data[971] = 8'b11111111;
  assign alpha_arctangen_expected_table_data[972] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[973] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[974] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[975] = 8'b00000001;
  assign alpha_arctangen_expected_table_data[976] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[977] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[978] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[979] = 8'b00000000;
  assign alpha_arctangen_expected_table_data[980] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[981] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[982] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[983] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[984] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[985] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[986] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[987] = 8'b00110010;
  assign alpha_arctangen_expected_table_data[988] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[989] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[990] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[991] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[992] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[993] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[994] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[995] = 8'b00110011;
  assign alpha_arctangen_expected_table_data[996] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[997] = 8'b01100100;
  assign alpha_arctangen_expected_table_data[998] = 8'b10011011;
  assign alpha_arctangen_expected_table_data[999] = 8'b10011100;
  assign alpha_arctangen_expected_table_data[1000] = 8'b10011100;
  assign alpha_arctangen_expected_1 = alpha_arctangen_expected_table_data[magnitude_addr];



  assign alpha_arctangen_expected_2 = alpha_arctangen_expected_1;



  assign alpha_arctangen_ref = alpha_arctangen_expected_2;

  always @(posedge clk)
    begin : alpha_arctangen_checker
      if (reset_x == 1'b1) begin
        alpha_arctangen_testFailure <= 1'b0;
      end
      else begin
        if (clk_enable == 1'b1 && alpha_arctangen !== alpha_arctangen_ref) begin
          alpha_arctangen_testFailure <= 1'b1;
          $display("ERROR in alpha_arctangen at time %t : Expected '%h' Actual '%h'", $time, alpha_arctangen_ref, alpha_arctangen);
        end
      end
    end

  assign testFailure = magnitude_testFailure | alpha_arctangen_testFailure;



  always @(posedge clk)
    begin : completed_msg
      if (snkDone == 1'b1) begin
        if (testFailure == 1'b0) begin
          $display("**************TEST COMPLETED (PASSED)**************");
        end
        else begin
          $display("**************TEST COMPLETED (FAILED)**************");
        end
      end
    end

endmodule  // simulink_functio_tb

